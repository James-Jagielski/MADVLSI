magic
tech sky130A
timestamp 1697759168
<< nwell >>
rect 770 2895 2670 2900
rect 370 2860 2670 2895
rect 350 2220 2690 2860
rect 370 2190 2670 2220
rect 445 2185 2670 2190
rect 745 2145 2670 2185
rect 750 2125 2670 2145
rect 900 2030 2670 2125
rect 900 1390 2690 2030
<< nmos >>
rect 870 645 920 1245
rect 970 645 1020 1245
rect 1070 645 1120 1245
rect 1170 645 1220 1245
rect 1270 645 1320 1245
rect 1345 645 1395 1245
rect 1420 645 1470 1245
rect 1495 645 1545 1245
rect 1570 645 1620 1245
rect 1645 645 1695 1245
rect 1745 645 1795 1245
rect 1820 645 1870 1245
rect 1895 645 1945 1245
rect 1970 645 2020 1245
rect 2045 645 2095 1245
rect 2120 645 2170 1245
rect 2220 645 2270 1245
rect 2320 645 2370 1245
rect 2420 645 2470 1245
rect 2520 645 2570 1245
rect 1020 -130 1070 470
rect 1120 -130 1170 470
rect 1220 -130 1270 470
rect 1320 -130 1370 470
rect 1420 -130 1470 470
rect 1520 -130 1570 470
rect 1620 -130 1670 470
rect 1720 -130 1770 470
rect 1820 -130 1870 470
rect 1920 -130 1970 470
rect 2020 -130 2070 470
rect 2120 -130 2170 470
rect 2220 -130 2270 470
rect 2320 -130 2370 470
rect 2420 -130 2470 470
rect 2520 -130 2570 470
<< pmos >>
rect 470 2240 520 2840
rect 570 2240 620 2840
rect 670 2240 720 2840
rect 770 2240 820 2840
rect 870 2240 920 2840
rect 970 2240 1020 2840
rect 1070 2240 1120 2840
rect 1145 2240 1195 2840
rect 1220 2240 1270 2840
rect 1295 2240 1345 2840
rect 1370 2240 1420 2840
rect 1445 2240 1495 2840
rect 1545 2240 1595 2840
rect 1620 2240 1670 2840
rect 1695 2240 1745 2840
rect 1770 2240 1820 2840
rect 1845 2240 1895 2840
rect 1920 2240 1970 2840
rect 2020 2240 2070 2840
rect 2120 2240 2170 2840
rect 2220 2240 2270 2840
rect 2320 2240 2370 2840
rect 2420 2240 2470 2840
rect 2520 2240 2570 2840
rect 1020 1410 1070 2010
rect 1120 1410 1170 2010
rect 1220 1410 1270 2010
rect 1320 1410 1370 2010
rect 1420 1410 1470 2010
rect 1520 1410 1570 2010
rect 1620 1410 1670 2010
rect 1720 1410 1770 2010
rect 1820 1410 1870 2010
rect 1920 1410 1970 2010
rect 2020 1410 2070 2010
rect 2120 1410 2170 2010
rect 2220 1410 2270 2010
rect 2320 1410 2370 2010
rect 2420 1410 2470 2010
rect 2520 1410 2570 2010
<< ndiff >>
rect 820 1235 870 1245
rect 820 660 835 1235
rect 855 660 870 1235
rect 820 645 870 660
rect 920 1235 970 1245
rect 920 660 935 1235
rect 955 660 970 1235
rect 920 645 970 660
rect 1020 1235 1070 1245
rect 1020 660 1035 1235
rect 1055 660 1070 1235
rect 1020 645 1070 660
rect 1120 1235 1170 1245
rect 1120 660 1135 1235
rect 1155 660 1170 1235
rect 1120 645 1170 660
rect 1220 1235 1270 1245
rect 1220 660 1235 1235
rect 1255 660 1270 1235
rect 1220 645 1270 660
rect 1320 645 1345 1245
rect 1395 645 1420 1245
rect 1470 645 1495 1245
rect 1545 645 1570 1245
rect 1620 645 1645 1245
rect 1695 1235 1745 1245
rect 1695 660 1710 1235
rect 1730 660 1745 1235
rect 1695 645 1745 660
rect 1795 645 1820 1245
rect 1870 645 1895 1245
rect 1945 645 1970 1245
rect 2020 645 2045 1245
rect 2095 645 2120 1245
rect 2170 1235 2220 1245
rect 2170 660 2185 1235
rect 2205 660 2220 1235
rect 2170 645 2220 660
rect 2270 1235 2320 1245
rect 2270 660 2285 1235
rect 2305 660 2320 1235
rect 2270 645 2320 660
rect 2370 1235 2420 1245
rect 2370 660 2385 1235
rect 2405 660 2420 1235
rect 2370 645 2420 660
rect 2470 1235 2520 1245
rect 2470 660 2485 1235
rect 2505 660 2520 1235
rect 2470 645 2520 660
rect 2570 1235 2620 1245
rect 2570 660 2585 1235
rect 2605 660 2620 1235
rect 2570 645 2620 660
rect 970 460 1020 470
rect 970 -115 985 460
rect 1005 -115 1020 460
rect 970 -130 1020 -115
rect 1070 460 1120 470
rect 1070 -115 1085 460
rect 1105 -115 1120 460
rect 1070 -130 1120 -115
rect 1170 460 1220 470
rect 1170 -115 1185 460
rect 1205 -115 1220 460
rect 1170 -130 1220 -115
rect 1270 460 1320 470
rect 1270 -115 1285 460
rect 1305 -115 1320 460
rect 1270 -130 1320 -115
rect 1370 460 1420 470
rect 1370 -115 1385 460
rect 1405 -115 1420 460
rect 1370 -130 1420 -115
rect 1470 460 1520 470
rect 1470 -115 1485 460
rect 1505 -115 1520 460
rect 1470 -130 1520 -115
rect 1570 460 1620 470
rect 1570 -115 1585 460
rect 1605 -115 1620 460
rect 1570 -130 1620 -115
rect 1670 460 1720 470
rect 1670 -115 1685 460
rect 1705 -115 1720 460
rect 1670 -130 1720 -115
rect 1770 460 1820 470
rect 1770 -115 1785 460
rect 1805 -115 1820 460
rect 1770 -130 1820 -115
rect 1870 460 1920 470
rect 1870 -115 1885 460
rect 1905 -115 1920 460
rect 1870 -130 1920 -115
rect 1970 460 2020 470
rect 1970 -115 1985 460
rect 2005 -115 2020 460
rect 1970 -130 2020 -115
rect 2070 460 2120 470
rect 2070 -115 2085 460
rect 2105 -115 2120 460
rect 2070 -130 2120 -115
rect 2170 460 2220 470
rect 2170 -115 2185 460
rect 2205 -115 2220 460
rect 2170 -130 2220 -115
rect 2270 460 2320 470
rect 2270 -115 2285 460
rect 2305 -115 2320 460
rect 2270 -130 2320 -115
rect 2370 460 2420 470
rect 2370 -115 2385 460
rect 2405 -115 2420 460
rect 2370 -130 2420 -115
rect 2470 460 2520 470
rect 2470 -115 2485 460
rect 2505 -115 2520 460
rect 2470 -130 2520 -115
rect 2570 460 2620 470
rect 2570 -115 2585 460
rect 2605 -115 2620 460
rect 2570 -130 2620 -115
<< pdiff >>
rect 420 2830 470 2840
rect 420 2255 435 2830
rect 455 2255 470 2830
rect 420 2240 470 2255
rect 520 2830 570 2840
rect 520 2255 535 2830
rect 555 2255 570 2830
rect 520 2240 570 2255
rect 620 2830 670 2840
rect 620 2255 635 2830
rect 655 2255 670 2830
rect 620 2240 670 2255
rect 720 2830 770 2840
rect 720 2255 735 2830
rect 755 2255 770 2830
rect 720 2240 770 2255
rect 820 2830 870 2840
rect 820 2255 835 2830
rect 855 2255 870 2830
rect 820 2240 870 2255
rect 920 2830 970 2840
rect 920 2255 935 2830
rect 955 2255 970 2830
rect 920 2240 970 2255
rect 1020 2830 1070 2840
rect 1020 2255 1035 2830
rect 1055 2255 1070 2830
rect 1020 2240 1070 2255
rect 1120 2240 1145 2840
rect 1195 2240 1220 2840
rect 1270 2240 1295 2840
rect 1345 2240 1370 2840
rect 1420 2240 1445 2840
rect 1495 2825 1545 2840
rect 1495 2255 1510 2825
rect 1530 2255 1545 2825
rect 1495 2240 1545 2255
rect 1595 2240 1620 2840
rect 1670 2240 1695 2840
rect 1745 2240 1770 2840
rect 1820 2240 1845 2840
rect 1895 2240 1920 2840
rect 1970 2830 2020 2840
rect 1970 2255 1985 2830
rect 2005 2255 2020 2830
rect 1970 2240 2020 2255
rect 2070 2830 2120 2840
rect 2070 2255 2085 2830
rect 2105 2255 2120 2830
rect 2070 2240 2120 2255
rect 2170 2830 2220 2840
rect 2170 2255 2185 2830
rect 2205 2255 2220 2830
rect 2170 2240 2220 2255
rect 2270 2830 2320 2840
rect 2270 2255 2285 2830
rect 2305 2255 2320 2830
rect 2270 2240 2320 2255
rect 2370 2830 2420 2840
rect 2370 2255 2385 2830
rect 2405 2255 2420 2830
rect 2370 2240 2420 2255
rect 2470 2830 2520 2840
rect 2470 2255 2485 2830
rect 2505 2255 2520 2830
rect 2470 2240 2520 2255
rect 2570 2830 2620 2840
rect 2570 2255 2585 2830
rect 2605 2255 2620 2830
rect 2570 2240 2620 2255
rect 970 2000 1020 2010
rect 970 1425 985 2000
rect 1005 1425 1020 2000
rect 970 1410 1020 1425
rect 1070 2000 1120 2010
rect 1070 1425 1085 2000
rect 1105 1425 1120 2000
rect 1070 1410 1120 1425
rect 1170 2000 1220 2010
rect 1170 1425 1185 2000
rect 1205 1425 1220 2000
rect 1170 1410 1220 1425
rect 1270 2000 1320 2010
rect 1270 1425 1285 2000
rect 1305 1425 1320 2000
rect 1270 1410 1320 1425
rect 1370 2000 1420 2010
rect 1370 1425 1385 2000
rect 1405 1425 1420 2000
rect 1370 1410 1420 1425
rect 1470 2000 1520 2010
rect 1470 1425 1485 2000
rect 1505 1425 1520 2000
rect 1470 1410 1520 1425
rect 1570 2000 1620 2010
rect 1570 1425 1585 2000
rect 1605 1425 1620 2000
rect 1570 1410 1620 1425
rect 1670 2000 1720 2010
rect 1670 1425 1685 2000
rect 1705 1425 1720 2000
rect 1670 1410 1720 1425
rect 1770 2000 1820 2010
rect 1770 1425 1785 2000
rect 1805 1425 1820 2000
rect 1770 1410 1820 1425
rect 1870 2000 1920 2010
rect 1870 1425 1885 2000
rect 1905 1425 1920 2000
rect 1870 1410 1920 1425
rect 1970 2000 2020 2010
rect 1970 1425 1985 2000
rect 2005 1425 2020 2000
rect 1970 1410 2020 1425
rect 2070 2000 2120 2010
rect 2070 1425 2085 2000
rect 2105 1425 2120 2000
rect 2070 1410 2120 1425
rect 2170 2000 2220 2010
rect 2170 1425 2185 2000
rect 2205 1425 2220 2000
rect 2170 1410 2220 1425
rect 2270 2000 2320 2010
rect 2270 1425 2285 2000
rect 2305 1425 2320 2000
rect 2270 1410 2320 1425
rect 2370 2000 2420 2010
rect 2370 1425 2385 2000
rect 2405 1425 2420 2000
rect 2370 1410 2420 1425
rect 2470 2000 2520 2010
rect 2470 1425 2485 2000
rect 2505 1425 2520 2000
rect 2470 1410 2520 1425
rect 2570 2000 2620 2010
rect 2570 1425 2585 2000
rect 2605 1425 2620 2000
rect 2570 1410 2620 1425
<< ndiffc >>
rect 835 660 855 1235
rect 935 660 955 1235
rect 1035 660 1055 1235
rect 1135 660 1155 1235
rect 1235 660 1255 1235
rect 1710 660 1730 1235
rect 2185 660 2205 1235
rect 2285 660 2305 1235
rect 2385 660 2405 1235
rect 2485 660 2505 1235
rect 2585 660 2605 1235
rect 985 -115 1005 460
rect 1085 -115 1105 460
rect 1185 -115 1205 460
rect 1285 -115 1305 460
rect 1385 -115 1405 460
rect 1485 -115 1505 460
rect 1585 -115 1605 460
rect 1685 -115 1705 460
rect 1785 -115 1805 460
rect 1885 -115 1905 460
rect 1985 -115 2005 460
rect 2085 -115 2105 460
rect 2185 -115 2205 460
rect 2285 -115 2305 460
rect 2385 -115 2405 460
rect 2485 -115 2505 460
rect 2585 -115 2605 460
<< pdiffc >>
rect 435 2255 455 2830
rect 535 2255 555 2830
rect 635 2255 655 2830
rect 735 2255 755 2830
rect 835 2255 855 2830
rect 935 2255 955 2830
rect 1035 2255 1055 2830
rect 1510 2255 1530 2825
rect 1985 2255 2005 2830
rect 2085 2255 2105 2830
rect 2185 2255 2205 2830
rect 2285 2255 2305 2830
rect 2385 2255 2405 2830
rect 2485 2255 2505 2830
rect 2585 2255 2605 2830
rect 985 1425 1005 2000
rect 1085 1425 1105 2000
rect 1185 1425 1205 2000
rect 1285 1425 1305 2000
rect 1385 1425 1405 2000
rect 1485 1425 1505 2000
rect 1585 1425 1605 2000
rect 1685 1425 1705 2000
rect 1785 1425 1805 2000
rect 1885 1425 1905 2000
rect 1985 1425 2005 2000
rect 2085 1425 2105 2000
rect 2185 1425 2205 2000
rect 2285 1425 2305 2000
rect 2385 1425 2405 2000
rect 2485 1425 2505 2000
rect 2585 1425 2605 2000
<< psubdiff >>
rect 770 1235 820 1245
rect 770 660 785 1235
rect 805 660 820 1235
rect 770 645 820 660
rect 2620 1235 2670 1245
rect 2620 660 2635 1235
rect 2655 660 2670 1235
rect 2620 645 2670 660
rect 920 460 970 470
rect 920 -115 935 460
rect 955 -115 970 460
rect 920 -130 970 -115
rect 2620 460 2670 470
rect 2620 -115 2635 460
rect 2655 -115 2670 460
rect 2620 -130 2670 -115
<< nsubdiff >>
rect 370 2830 420 2840
rect 370 2255 385 2830
rect 405 2255 420 2830
rect 370 2240 420 2255
rect 2620 2830 2670 2840
rect 2620 2255 2635 2830
rect 2655 2255 2670 2830
rect 2620 2240 2670 2255
rect 920 2000 970 2010
rect 920 1425 935 2000
rect 955 1425 970 2000
rect 920 1410 970 1425
rect 2620 2000 2670 2010
rect 2620 1425 2635 2000
rect 2655 1425 2670 2000
rect 2620 1410 2670 1425
<< psubdiffcont >>
rect 785 660 805 1235
rect 2635 660 2655 1235
rect 935 -115 955 460
rect 2635 -115 2655 460
<< nsubdiffcont >>
rect 385 2255 405 2830
rect 2635 2255 2655 2830
rect 935 1425 955 2000
rect 2635 1425 2655 2000
<< poly >>
rect 475 2885 515 2895
rect 475 2865 485 2885
rect 505 2865 515 2885
rect 475 2855 515 2865
rect 545 2885 2495 2895
rect 545 2865 555 2885
rect 575 2880 2465 2885
rect 575 2865 620 2880
rect 545 2855 620 2865
rect 470 2840 520 2855
rect 570 2840 620 2855
rect 670 2840 720 2880
rect 770 2840 820 2855
rect 870 2840 920 2880
rect 970 2840 1020 2855
rect 1070 2840 1120 2880
rect 1145 2840 1195 2880
rect 1220 2840 1270 2880
rect 1295 2840 1345 2880
rect 1370 2840 1420 2880
rect 1445 2840 1495 2880
rect 1545 2840 1595 2880
rect 1620 2840 1670 2880
rect 1695 2840 1745 2880
rect 1770 2840 1820 2880
rect 1845 2840 1895 2880
rect 1920 2840 1970 2880
rect 2020 2840 2070 2855
rect 2120 2840 2170 2880
rect 2220 2840 2270 2855
rect 2320 2840 2370 2880
rect 2420 2865 2465 2880
rect 2485 2865 2495 2885
rect 2420 2855 2495 2865
rect 2525 2885 2565 2895
rect 2525 2865 2535 2885
rect 2555 2865 2565 2885
rect 2525 2855 2565 2865
rect 2420 2840 2470 2855
rect 2520 2840 2570 2855
rect 470 2225 520 2240
rect 570 2225 620 2240
rect 670 2225 720 2240
rect 770 2225 820 2240
rect 870 2225 920 2240
rect 970 2225 1020 2240
rect 1070 2225 1120 2240
rect 1145 2225 1195 2240
rect 1220 2225 1270 2240
rect 1295 2225 1345 2240
rect 1370 2225 1420 2240
rect 1445 2225 1495 2240
rect 1545 2225 1595 2240
rect 1620 2225 1670 2240
rect 1695 2225 1745 2240
rect 1770 2225 1820 2240
rect 1845 2225 1895 2240
rect 1920 2225 1970 2240
rect 2020 2225 2070 2240
rect 2120 2225 2170 2240
rect 2220 2225 2270 2240
rect 2320 2225 2370 2240
rect 2420 2225 2470 2240
rect 2520 2225 2570 2240
rect 775 2215 815 2225
rect 775 2195 785 2215
rect 805 2195 815 2215
rect 775 2185 815 2195
rect 980 2215 1020 2225
rect 980 2195 990 2215
rect 1010 2195 1020 2215
rect 980 2185 1020 2195
rect 2025 2215 2065 2225
rect 2025 2195 2035 2215
rect 2055 2195 2065 2215
rect 2025 2185 2065 2195
rect 2225 2215 2265 2225
rect 2225 2195 2235 2215
rect 2255 2195 2265 2215
rect 2225 2185 2265 2195
rect 1120 2105 2460 2120
rect 1120 2065 1135 2105
rect 2445 2065 2460 2105
rect 995 2055 1035 2065
rect 995 2035 1005 2055
rect 1025 2035 1035 2055
rect 675 2025 715 2035
rect 995 2025 1035 2035
rect 1095 2055 1135 2065
rect 1095 2035 1105 2055
rect 1125 2035 1135 2055
rect 1095 2025 1135 2035
rect 1255 2055 1295 2065
rect 1255 2035 1265 2055
rect 1285 2035 1295 2055
rect 1475 2055 1515 2065
rect 1475 2040 1485 2055
rect 1255 2025 1295 2035
rect 1320 2035 1485 2040
rect 1505 2040 1515 2055
rect 1675 2055 1715 2065
rect 1675 2040 1685 2055
rect 1505 2035 1685 2040
rect 1705 2040 1715 2055
rect 1875 2055 1915 2065
rect 1875 2040 1885 2055
rect 1705 2035 1885 2040
rect 1905 2040 1915 2055
rect 2075 2055 2115 2065
rect 2075 2040 2085 2055
rect 1905 2035 2085 2040
rect 2105 2040 2115 2055
rect 2295 2055 2335 2065
rect 2105 2035 2270 2040
rect 1320 2025 2270 2035
rect 2295 2035 2305 2055
rect 2325 2035 2335 2055
rect 2295 2025 2335 2035
rect 2430 2055 2470 2065
rect 2430 2035 2440 2055
rect 2460 2035 2470 2055
rect 2430 2025 2470 2035
rect 2555 2055 2595 2065
rect 2555 2035 2565 2055
rect 2585 2035 2595 2055
rect 2555 2025 2595 2035
rect 675 2005 685 2025
rect 705 2005 715 2025
rect 1020 2010 1070 2025
rect 1120 2010 1170 2025
rect 1220 2010 1270 2025
rect 1320 2010 1370 2025
rect 1420 2010 1470 2025
rect 1520 2010 1570 2025
rect 1620 2010 1670 2025
rect 1720 2010 1770 2025
rect 1820 2010 1870 2025
rect 1920 2010 1970 2025
rect 2020 2010 2070 2025
rect 2120 2010 2170 2025
rect 2220 2010 2270 2025
rect 2320 2010 2370 2025
rect 2420 2010 2470 2025
rect 2520 2010 2570 2025
rect 675 1995 715 2005
rect 700 1345 715 1995
rect 1020 1395 1070 1410
rect 1120 1395 1170 1410
rect 1220 1395 1270 1410
rect 1320 1395 1370 1410
rect 1420 1395 1470 1410
rect 1520 1395 1570 1410
rect 1620 1395 1670 1410
rect 1720 1395 1770 1410
rect 1820 1395 1870 1410
rect 1920 1395 1970 1410
rect 2020 1395 2070 1410
rect 2120 1395 2170 1410
rect 2220 1395 2270 1410
rect 2320 1395 2370 1410
rect 2420 1395 2470 1410
rect 2520 1395 2570 1410
rect 1535 1350 1550 1395
rect 695 1330 960 1345
rect 1535 1340 1740 1350
rect 1535 1335 1710 1340
rect 945 1300 960 1330
rect 1700 1320 1710 1335
rect 1730 1320 1740 1340
rect 1700 1310 1740 1320
rect 845 1290 885 1300
rect 845 1270 855 1290
rect 875 1270 885 1290
rect 845 1260 885 1270
rect 945 1290 1680 1300
rect 945 1270 955 1290
rect 975 1285 1680 1290
rect 1760 1290 2495 1300
rect 1760 1285 2465 1290
rect 975 1270 1020 1285
rect 945 1260 1020 1270
rect 870 1245 920 1260
rect 970 1245 1020 1260
rect 1070 1245 1120 1285
rect 1170 1245 1220 1260
rect 1270 1245 1320 1285
rect 1345 1245 1395 1285
rect 1420 1245 1470 1285
rect 1495 1245 1545 1285
rect 1570 1245 1620 1285
rect 1645 1270 1795 1285
rect 1645 1245 1695 1270
rect 1745 1245 1795 1270
rect 1820 1245 1870 1285
rect 1895 1245 1945 1285
rect 1970 1245 2020 1285
rect 2045 1245 2095 1285
rect 2120 1245 2170 1285
rect 2220 1245 2270 1260
rect 2320 1245 2370 1285
rect 2420 1270 2465 1285
rect 2485 1270 2495 1290
rect 2420 1260 2495 1270
rect 2555 1290 2595 1300
rect 2555 1270 2565 1290
rect 2585 1270 2595 1290
rect 2555 1260 2595 1270
rect 2420 1245 2470 1260
rect 2520 1245 2570 1260
rect 870 630 920 645
rect 970 630 1020 645
rect 1070 630 1120 645
rect 1170 630 1220 645
rect 1270 630 1320 645
rect 1345 630 1395 645
rect 1420 630 1470 645
rect 1495 630 1545 645
rect 1570 630 1620 645
rect 1645 630 1695 645
rect 1745 630 1795 645
rect 1820 630 1870 645
rect 1895 630 1945 645
rect 1970 630 2020 645
rect 2045 630 2095 645
rect 2120 630 2170 645
rect 2220 630 2270 645
rect 2320 630 2370 645
rect 2420 630 2470 645
rect 2520 630 2570 645
rect 1170 620 1210 630
rect 1170 600 1180 620
rect 1200 600 1210 620
rect 1170 590 1210 600
rect 2195 620 2235 630
rect 2195 600 2205 620
rect 2225 600 2235 620
rect 2195 590 2235 600
rect 995 515 1035 525
rect 995 495 1005 515
rect 1025 495 1035 515
rect 995 485 1035 495
rect 1095 515 1135 525
rect 1095 495 1105 515
rect 1125 495 1135 515
rect 1095 485 1135 495
rect 1255 515 1295 525
rect 1255 495 1265 515
rect 1285 495 1295 515
rect 1475 515 1515 525
rect 1475 500 1485 515
rect 1255 485 1295 495
rect 1320 495 1485 500
rect 1505 500 1515 515
rect 1675 515 1715 525
rect 1675 500 1685 515
rect 1505 495 1685 500
rect 1705 500 1715 515
rect 1875 515 1915 525
rect 1875 500 1885 515
rect 1705 495 1885 500
rect 1905 500 1915 515
rect 2075 515 2115 525
rect 2075 500 2085 515
rect 1905 495 2085 500
rect 2105 500 2115 515
rect 2295 515 2335 525
rect 2105 495 2270 500
rect 1320 485 2270 495
rect 2295 495 2305 515
rect 2325 495 2335 515
rect 2295 485 2335 495
rect 2425 515 2465 530
rect 2425 495 2435 515
rect 2455 495 2465 515
rect 2425 485 2465 495
rect 2555 515 2595 525
rect 2555 495 2565 515
rect 2585 495 2595 515
rect 2555 485 2595 495
rect 1020 470 1070 485
rect 1120 470 1170 485
rect 1220 470 1270 485
rect 1320 470 1370 485
rect 1420 470 1470 485
rect 1520 470 1570 485
rect 1620 470 1670 485
rect 1720 470 1770 485
rect 1820 470 1870 485
rect 1920 470 1970 485
rect 2020 470 2070 485
rect 2120 470 2170 485
rect 2220 470 2270 485
rect 2320 470 2370 485
rect 2420 470 2470 485
rect 2520 470 2570 485
rect 1020 -145 1070 -130
rect 1120 -145 1170 -130
rect 1220 -145 1270 -130
rect 1320 -145 1370 -130
rect 1420 -145 1470 -130
rect 1520 -145 1570 -130
rect 1620 -145 1670 -130
rect 1720 -145 1770 -130
rect 1820 -145 1870 -130
rect 1920 -145 1970 -130
rect 2020 -145 2070 -130
rect 2120 -145 2170 -130
rect 2220 -145 2270 -130
rect 2320 -145 2370 -130
rect 2420 -145 2470 -130
rect 2520 -145 2570 -130
<< polycont >>
rect 485 2865 505 2885
rect 555 2865 575 2885
rect 2465 2865 2485 2885
rect 2535 2865 2555 2885
rect 785 2195 805 2215
rect 990 2195 1010 2215
rect 2035 2195 2055 2215
rect 2235 2195 2255 2215
rect 1005 2035 1025 2055
rect 1105 2035 1125 2055
rect 1265 2035 1285 2055
rect 1485 2035 1505 2055
rect 1685 2035 1705 2055
rect 1885 2035 1905 2055
rect 2085 2035 2105 2055
rect 2305 2035 2325 2055
rect 2440 2035 2460 2055
rect 2565 2035 2585 2055
rect 685 2005 705 2025
rect 1710 1320 1730 1340
rect 855 1270 875 1290
rect 955 1270 975 1290
rect 2465 1270 2485 1290
rect 2565 1270 2585 1290
rect 1180 600 1200 620
rect 2205 600 2225 620
rect 1005 495 1025 515
rect 1105 495 1125 515
rect 1265 495 1285 515
rect 1485 495 1505 515
rect 1685 495 1705 515
rect 1885 495 1905 515
rect 2085 495 2105 515
rect 2305 495 2325 515
rect 2435 495 2455 515
rect 2565 495 2585 515
<< locali >>
rect 745 2910 2305 2930
rect 475 2885 515 2895
rect 475 2875 485 2885
rect 445 2865 485 2875
rect 505 2865 515 2885
rect 445 2855 515 2865
rect 545 2885 585 2895
rect 545 2865 555 2885
rect 575 2865 585 2885
rect 545 2855 585 2865
rect 445 2835 465 2855
rect 545 2835 565 2855
rect 745 2835 765 2910
rect 945 2855 2105 2875
rect 945 2835 965 2855
rect 2085 2835 2105 2855
rect 2285 2835 2305 2910
rect 2455 2885 2495 2895
rect 2455 2865 2465 2885
rect 2485 2865 2495 2885
rect 2455 2855 2495 2865
rect 2525 2885 2565 2895
rect 2525 2865 2535 2885
rect 2555 2875 2565 2885
rect 2555 2865 2595 2875
rect 2525 2855 2595 2865
rect 2475 2835 2495 2855
rect 2575 2835 2595 2855
rect 375 2830 465 2835
rect 375 2255 385 2830
rect 405 2255 435 2830
rect 455 2255 465 2830
rect 375 2245 465 2255
rect 525 2830 565 2835
rect 525 2255 535 2830
rect 555 2255 565 2830
rect 525 2245 565 2255
rect 625 2830 665 2835
rect 625 2255 635 2830
rect 655 2255 665 2830
rect 625 2245 665 2255
rect 725 2830 765 2835
rect 725 2255 735 2830
rect 755 2255 765 2830
rect 725 2245 765 2255
rect 825 2830 865 2835
rect 825 2255 835 2830
rect 855 2255 865 2830
rect 825 2245 865 2255
rect 925 2830 965 2835
rect 925 2255 935 2830
rect 955 2255 965 2830
rect 925 2245 965 2255
rect 1025 2830 1065 2835
rect 1025 2255 1035 2830
rect 1055 2255 1065 2830
rect 1025 2245 1065 2255
rect 1500 2825 1540 2835
rect 1500 2255 1510 2825
rect 1530 2255 1540 2825
rect 1500 2245 1540 2255
rect 1975 2830 2015 2835
rect 1975 2255 1985 2830
rect 2005 2255 2015 2830
rect 1975 2245 2015 2255
rect 2075 2830 2115 2835
rect 2075 2255 2085 2830
rect 2105 2255 2115 2830
rect 2075 2245 2115 2255
rect 2175 2830 2215 2835
rect 2175 2255 2185 2830
rect 2205 2255 2215 2830
rect 2175 2245 2215 2255
rect 2275 2830 2315 2835
rect 2275 2255 2285 2830
rect 2305 2255 2315 2830
rect 2275 2245 2315 2255
rect 2375 2830 2415 2835
rect 2375 2255 2385 2830
rect 2405 2255 2415 2830
rect 2375 2245 2415 2255
rect 2475 2830 2515 2835
rect 2475 2255 2485 2830
rect 2505 2255 2515 2830
rect 2475 2245 2515 2255
rect 2575 2830 2665 2835
rect 2575 2255 2585 2830
rect 2605 2255 2635 2830
rect 2655 2255 2665 2830
rect 2575 2245 2665 2255
rect 535 2175 555 2245
rect 725 2220 745 2245
rect 825 2225 845 2245
rect 350 2155 555 2175
rect 680 2200 745 2220
rect 775 2215 845 2225
rect 680 2035 700 2200
rect 775 2195 785 2215
rect 805 2205 845 2215
rect 805 2195 815 2205
rect 775 2185 815 2195
rect 925 2165 945 2245
rect 1030 2225 1050 2245
rect 980 2215 1050 2225
rect 980 2195 990 2215
rect 1010 2205 1050 2215
rect 1010 2195 1020 2205
rect 980 2185 1020 2195
rect 1500 2180 1520 2245
rect 1990 2225 2010 2245
rect 2190 2225 2210 2245
rect 1990 2215 2065 2225
rect 1990 2205 2035 2215
rect 2025 2195 2035 2205
rect 2055 2195 2065 2215
rect 2190 2215 2265 2225
rect 2190 2205 2235 2215
rect 2025 2185 2065 2195
rect 2225 2195 2235 2205
rect 2255 2195 2265 2215
rect 2225 2185 2265 2195
rect 735 2145 945 2165
rect 1040 2160 1520 2180
rect 2490 2175 2510 2245
rect 675 2025 715 2035
rect 675 2005 685 2025
rect 705 2005 715 2025
rect 675 1995 715 2005
rect 735 1975 755 2145
rect 1040 2115 1060 2160
rect 2490 2155 2725 2175
rect 695 1950 755 1975
rect 780 2095 1060 2115
rect 695 -160 715 1950
rect 780 1325 800 2095
rect 1185 2085 2405 2105
rect 995 2055 1035 2065
rect 995 2035 1005 2055
rect 1025 2035 1035 2055
rect 995 2025 1035 2035
rect 1095 2055 1135 2065
rect 1095 2035 1105 2055
rect 1125 2035 1135 2055
rect 1095 2025 1135 2035
rect 995 2005 1015 2025
rect 1095 2005 1115 2025
rect 1185 2005 1205 2085
rect 1255 2055 1295 2065
rect 1255 2035 1265 2055
rect 1285 2035 1295 2055
rect 1255 2025 1295 2035
rect 1275 2005 1295 2025
rect 1385 2005 1405 2085
rect 1475 2055 1515 2065
rect 1475 2035 1485 2055
rect 1505 2035 1515 2055
rect 1475 2025 1515 2035
rect 1485 2005 1505 2025
rect 1585 2005 1605 2085
rect 1675 2055 1715 2065
rect 1675 2035 1685 2055
rect 1705 2035 1715 2055
rect 1675 2025 1715 2035
rect 1685 2005 1705 2025
rect 1785 2005 1805 2085
rect 1875 2055 1915 2065
rect 1875 2035 1885 2055
rect 1905 2035 1915 2055
rect 1875 2025 1915 2035
rect 1885 2005 1905 2025
rect 1985 2005 2005 2085
rect 2075 2055 2115 2065
rect 2075 2035 2085 2055
rect 2105 2035 2115 2055
rect 2075 2025 2115 2035
rect 2085 2005 2105 2025
rect 2185 2005 2205 2085
rect 2295 2055 2335 2065
rect 2295 2035 2305 2055
rect 2325 2035 2335 2055
rect 2295 2025 2335 2035
rect 2295 2005 2315 2025
rect 2385 2005 2405 2085
rect 2445 2085 2725 2105
rect 2445 2065 2465 2085
rect 2430 2055 2470 2065
rect 2430 2035 2440 2055
rect 2460 2045 2470 2055
rect 2555 2055 2595 2065
rect 2460 2035 2505 2045
rect 2430 2025 2505 2035
rect 2555 2035 2565 2055
rect 2585 2035 2595 2055
rect 2555 2025 2595 2035
rect 2485 2005 2505 2025
rect 2575 2005 2595 2025
rect 925 2000 1015 2005
rect 925 1425 935 2000
rect 955 1425 985 2000
rect 1005 1425 1015 2000
rect 925 1415 1015 1425
rect 1075 2000 1115 2005
rect 1075 1425 1085 2000
rect 1105 1425 1115 2000
rect 1075 1415 1115 1425
rect 1175 2000 1215 2005
rect 1175 1425 1185 2000
rect 1205 1425 1215 2000
rect 1175 1415 1215 1425
rect 1275 2000 1315 2005
rect 1275 1425 1285 2000
rect 1305 1425 1315 2000
rect 1275 1415 1315 1425
rect 1375 2000 1415 2005
rect 1375 1425 1385 2000
rect 1405 1425 1415 2000
rect 1375 1415 1415 1425
rect 1475 2000 1515 2005
rect 1475 1425 1485 2000
rect 1505 1425 1515 2000
rect 1475 1415 1515 1425
rect 1575 2000 1615 2005
rect 1575 1425 1585 2000
rect 1605 1425 1615 2000
rect 1575 1415 1615 1425
rect 1675 2000 1715 2005
rect 1675 1425 1685 2000
rect 1705 1425 1715 2000
rect 1675 1415 1715 1425
rect 1775 2000 1815 2005
rect 1775 1425 1785 2000
rect 1805 1425 1815 2000
rect 1775 1415 1815 1425
rect 1875 2000 1915 2005
rect 1875 1425 1885 2000
rect 1905 1425 1915 2000
rect 1875 1415 1915 1425
rect 1975 2000 2015 2005
rect 1975 1425 1985 2000
rect 2005 1425 2015 2000
rect 1975 1415 2015 1425
rect 2075 2000 2115 2005
rect 2075 1425 2085 2000
rect 2105 1425 2115 2000
rect 2075 1415 2115 1425
rect 2175 2000 2215 2005
rect 2175 1425 2185 2000
rect 2205 1425 2215 2000
rect 2175 1415 2215 1425
rect 2275 2000 2315 2005
rect 2275 1425 2285 2000
rect 2305 1425 2315 2000
rect 2275 1415 2315 1425
rect 2375 2000 2415 2005
rect 2375 1425 2385 2000
rect 2405 1425 2415 2000
rect 2375 1415 2415 1425
rect 2475 2000 2515 2005
rect 2475 1425 2485 2000
rect 2505 1425 2515 2000
rect 2475 1415 2515 1425
rect 2575 2000 2665 2005
rect 2575 1425 2585 2000
rect 2605 1425 2635 2000
rect 2655 1425 2665 2000
rect 2575 1415 2665 1425
rect 1085 1390 1105 1415
rect 2490 1390 2510 1415
rect 1085 1370 2510 1390
rect 735 1305 800 1325
rect 735 565 755 1305
rect 845 1290 885 1300
rect 845 1270 855 1290
rect 875 1270 885 1290
rect 845 1260 885 1270
rect 945 1290 985 1300
rect 945 1270 955 1290
rect 975 1270 985 1290
rect 945 1260 985 1270
rect 845 1240 865 1260
rect 945 1240 965 1260
rect 1145 1240 1165 1370
rect 1700 1340 1740 1350
rect 1700 1320 1710 1340
rect 1730 1320 1740 1340
rect 1700 1310 1740 1320
rect 1710 1240 1730 1310
rect 2295 1240 2315 1370
rect 2475 1320 2805 1340
rect 2475 1300 2495 1320
rect 2455 1290 2495 1300
rect 2455 1270 2465 1290
rect 2485 1270 2495 1290
rect 2455 1260 2495 1270
rect 2555 1290 2595 1300
rect 2555 1270 2565 1290
rect 2585 1270 2595 1290
rect 2555 1260 2595 1270
rect 2475 1240 2495 1260
rect 2575 1240 2595 1260
rect 775 1235 865 1240
rect 775 660 785 1235
rect 805 660 835 1235
rect 855 660 865 1235
rect 775 650 865 660
rect 925 1235 965 1240
rect 925 660 935 1235
rect 955 660 965 1235
rect 925 650 965 660
rect 1025 1235 1065 1240
rect 1025 660 1035 1235
rect 1055 660 1065 1235
rect 1025 650 1065 660
rect 1125 1235 1165 1240
rect 1125 660 1135 1235
rect 1155 660 1165 1235
rect 1125 650 1165 660
rect 1225 1235 1265 1240
rect 1225 660 1235 1235
rect 1255 660 1265 1235
rect 1225 650 1265 660
rect 1700 1235 1740 1240
rect 1700 660 1710 1235
rect 1730 660 1740 1235
rect 1700 650 1740 660
rect 2175 1235 2215 1240
rect 2175 660 2185 1235
rect 2205 660 2215 1235
rect 2175 650 2215 660
rect 2275 1235 2315 1240
rect 2275 660 2285 1235
rect 2305 660 2315 1235
rect 2275 650 2315 660
rect 2375 1235 2415 1240
rect 2375 660 2385 1235
rect 2405 660 2415 1235
rect 2375 650 2415 660
rect 2475 1235 2515 1240
rect 2475 660 2485 1235
rect 2505 660 2515 1235
rect 2475 650 2515 660
rect 2575 1235 2665 1240
rect 2575 660 2585 1235
rect 2605 660 2635 1235
rect 2655 660 2665 1235
rect 2575 650 2665 660
rect 1025 645 1045 650
rect 1225 630 1245 650
rect 1170 620 1245 630
rect 1170 600 1180 620
rect 1200 610 1245 620
rect 2195 630 2215 650
rect 2195 620 2235 630
rect 1200 600 1210 610
rect 1170 590 1210 600
rect 2195 600 2205 620
rect 2225 600 2235 620
rect 2195 590 2235 600
rect 735 545 2100 565
rect 1475 525 1495 545
rect 2080 525 2100 545
rect 2445 550 2875 570
rect 2445 530 2465 550
rect 995 515 1035 525
rect 995 495 1005 515
rect 1025 495 1035 515
rect 995 485 1035 495
rect 1095 515 1135 525
rect 1095 495 1105 515
rect 1125 495 1135 515
rect 1095 485 1135 495
rect 1255 515 1295 525
rect 1255 495 1265 515
rect 1285 495 1295 515
rect 1255 485 1295 495
rect 1475 515 1515 525
rect 1475 495 1485 515
rect 1505 495 1515 515
rect 1475 485 1515 495
rect 1675 515 1715 525
rect 1675 495 1685 515
rect 1705 495 1715 515
rect 1675 485 1715 495
rect 1875 515 1915 525
rect 1875 495 1885 515
rect 1905 495 1915 515
rect 1875 485 1915 495
rect 2075 515 2115 525
rect 2075 495 2085 515
rect 2105 495 2115 515
rect 2075 485 2115 495
rect 2295 515 2335 525
rect 2295 495 2305 515
rect 2325 495 2335 515
rect 2295 485 2335 495
rect 2425 515 2465 530
rect 2555 515 2595 525
rect 2425 495 2435 515
rect 2455 495 2505 515
rect 2425 485 2465 495
rect 995 465 1015 485
rect 1095 465 1115 485
rect 1275 465 1295 485
rect 1485 465 1505 485
rect 1685 465 1705 485
rect 1885 465 1905 485
rect 2085 465 2105 485
rect 2295 465 2315 485
rect 2485 465 2505 495
rect 2555 495 2565 515
rect 2585 495 2595 515
rect 2555 485 2595 495
rect 2575 465 2595 485
rect 925 460 1015 465
rect 925 -115 935 460
rect 955 -115 985 460
rect 1005 -115 1015 460
rect 925 -125 1015 -115
rect 1075 460 1115 465
rect 1075 -115 1085 460
rect 1105 -115 1115 460
rect 1075 -125 1115 -115
rect 1175 460 1215 465
rect 1175 -115 1185 460
rect 1205 -115 1215 460
rect 1175 -125 1215 -115
rect 1275 460 1315 465
rect 1275 -115 1285 460
rect 1305 -115 1315 460
rect 1275 -125 1315 -115
rect 1375 460 1415 465
rect 1375 -115 1385 460
rect 1405 -115 1415 460
rect 1375 -125 1415 -115
rect 1475 460 1515 465
rect 1475 -115 1485 460
rect 1505 -115 1515 460
rect 1475 -125 1515 -115
rect 1575 460 1615 465
rect 1575 -115 1585 460
rect 1605 -115 1615 460
rect 1575 -125 1615 -115
rect 1675 460 1715 465
rect 1675 -115 1685 460
rect 1705 -115 1715 460
rect 1675 -125 1715 -115
rect 1775 460 1820 465
rect 1775 -115 1785 460
rect 1805 -115 1820 460
rect 1775 -125 1820 -115
rect 1875 460 1915 465
rect 1875 -115 1885 460
rect 1905 -115 1915 460
rect 1875 -125 1915 -115
rect 1975 460 2015 465
rect 1975 -115 1985 460
rect 2005 -115 2015 460
rect 1975 -125 2015 -115
rect 2075 460 2115 465
rect 2075 -115 2085 460
rect 2105 -115 2115 460
rect 2075 -125 2115 -115
rect 2175 460 2215 465
rect 2175 -115 2185 460
rect 2205 -115 2215 460
rect 2175 -125 2215 -115
rect 2275 460 2315 465
rect 2275 -115 2285 460
rect 2305 -115 2315 460
rect 2275 -125 2315 -115
rect 2375 460 2415 465
rect 2375 -115 2385 460
rect 2405 -115 2415 460
rect 2375 -125 2415 -115
rect 2475 460 2515 465
rect 2475 -115 2485 460
rect 2505 -115 2515 460
rect 2475 -125 2515 -115
rect 2575 460 2665 465
rect 2575 -115 2585 460
rect 2605 -115 2635 460
rect 2655 -115 2665 460
rect 2575 -125 2665 -115
rect 1080 -160 1105 -125
rect 695 -180 1105 -160
rect 1190 -145 1210 -125
rect 1385 -145 1405 -125
rect 1585 -145 1605 -125
rect 1785 -145 1805 -125
rect 1985 -145 2005 -125
rect 2185 -145 2205 -125
rect 2375 -145 2395 -125
rect 1190 -165 2395 -145
rect 1085 -185 1105 -180
rect 2485 -185 2505 -125
rect 1085 -205 2505 -185
<< viali >>
rect 385 2255 405 2830
rect 435 2255 455 2830
rect 635 2255 655 2830
rect 835 2255 855 2830
rect 1035 2255 1055 2830
rect 1985 2255 2005 2830
rect 2185 2255 2205 2830
rect 2385 2255 2405 2830
rect 2585 2255 2605 2830
rect 2635 2255 2655 2830
rect 935 1425 955 2000
rect 985 1425 1005 2000
rect 1285 1425 1305 2000
rect 2285 1425 2305 2000
rect 2585 1425 2605 2000
rect 2635 1425 2655 2000
rect 785 660 805 1235
rect 835 660 855 1235
rect 1035 660 1055 1235
rect 1235 660 1255 1235
rect 2185 660 2205 1235
rect 2385 660 2405 1235
rect 2585 660 2605 1235
rect 2635 660 2655 1235
rect 935 -115 955 460
rect 985 -115 1005 460
rect 1285 -115 1305 460
rect 2285 -115 2305 460
rect 2585 -115 2605 460
rect 2635 -115 2655 460
<< metal1 >>
rect 370 2835 2670 2840
rect 350 2830 2670 2835
rect 350 2255 385 2830
rect 405 2255 435 2830
rect 455 2255 635 2830
rect 655 2255 835 2830
rect 855 2255 1035 2830
rect 1055 2255 1985 2830
rect 2005 2255 2185 2830
rect 2205 2255 2385 2830
rect 2405 2255 2585 2830
rect 2605 2255 2635 2830
rect 2655 2255 2670 2830
rect 350 2245 2670 2255
rect 370 2240 2670 2245
rect 915 2000 2670 2010
rect 915 1425 935 2000
rect 955 1425 985 2000
rect 1005 1425 1285 2000
rect 1305 1425 2285 2000
rect 2305 1425 2585 2000
rect 2605 1425 2635 2000
rect 2655 1995 2670 2000
rect 2655 1695 2895 1995
rect 2655 1425 2670 1695
rect 915 1410 2670 1425
rect 725 1245 2670 1250
rect 375 1235 2670 1245
rect 375 660 785 1235
rect 805 660 835 1235
rect 855 660 1035 1235
rect 1055 660 1235 1235
rect 1255 660 2185 1235
rect 2205 660 2385 1235
rect 2405 660 2585 1235
rect 2605 660 2635 1235
rect 2655 905 2670 1235
rect 2655 660 2895 905
rect 375 605 2895 660
rect 375 590 2670 605
rect 755 580 2670 590
rect 765 460 2670 580
rect 765 -100 935 460
rect 780 -115 935 -100
rect 955 -115 985 460
rect 1005 -115 1285 460
rect 1305 -115 2285 460
rect 2305 -115 2585 460
rect 2605 -115 2635 460
rect 2655 -115 2670 460
rect 780 -135 2670 -115
<< labels >>
rlabel locali 2725 2165 2725 2165 3 Vbp
port 1 e
rlabel locali 2725 2095 2725 2095 3 Vcp
port 2 e
rlabel metal1 2895 1860 2895 1860 3 VDD
port 3 e
rlabel locali 2805 1330 2805 1330 3 Vbn
port 4 e
rlabel metal1 2895 765 2895 765 3 GND
port 5 e
rlabel locali 2875 560 2875 560 3 Vcn
port 6 e
<< end >>
