magic
tech sky130A
timestamp 1697759168
<< locali >>
rect -145 1610 20 1630
rect -180 1540 -100 1560
rect -120 1115 -100 1540
rect -5 1545 20 1610
rect -5 1525 70 1545
rect -120 1095 125 1115
rect -115 775 -20 795
rect -40 525 -20 775
rect -40 505 75 525
rect -95 5 130 25
use Cascode_voltage_bias  Cascode_voltage_bias_0
timestamp 1697759168
transform 1 0 -2825 0 1 -545
box 350 -205 2895 2930
use diffamp_cell  diffamp_cell_0
timestamp 1697759168
transform 1 0 95 0 1 1145
box -100 -1150 2040 400
<< end >>
