magic
tech sky130A
timestamp 1694484618
<< nwell >>
rect -125 135 85 375
<< nmos >>
rect -5 0 10 100
<< pmos >>
rect -5 155 10 355
<< ndiff >>
rect -55 85 -5 100
rect -55 15 -40 85
rect -20 15 -5 85
rect -55 0 -5 15
rect 10 85 60 100
rect 10 15 25 85
rect 45 15 60 85
rect 10 0 60 15
<< pdiff >>
rect -55 340 -5 355
rect -55 270 -40 340
rect -20 270 -5 340
rect -55 240 -5 270
rect -55 170 -40 240
rect -20 170 -5 240
rect -55 155 -5 170
rect 10 340 60 355
rect 10 270 25 340
rect 45 270 60 340
rect 10 240 60 270
rect 10 170 25 240
rect 45 170 60 240
rect 10 155 60 170
<< ndiffc >>
rect -40 15 -20 85
rect 25 15 45 85
<< pdiffc >>
rect -40 270 -20 340
rect -40 170 -20 240
rect 25 270 45 340
rect 25 170 45 240
<< psubdiff >>
rect -105 85 -55 100
rect -105 15 -90 85
rect -70 15 -55 85
rect -105 0 -55 15
<< nsubdiff >>
rect -105 340 -55 355
rect -105 270 -90 340
rect -70 270 -55 340
rect -105 240 -55 270
rect -105 170 -90 240
rect -70 170 -55 240
rect -105 155 -55 170
<< psubdiffcont >>
rect -90 15 -70 85
<< nsubdiffcont >>
rect -90 270 -70 340
rect -90 170 -70 240
<< poly >>
rect -5 355 10 370
rect -5 100 10 155
rect -5 -115 10 0
rect -30 -125 10 -115
rect -30 -145 -20 -125
rect 0 -145 10 -125
rect -30 -155 10 -145
<< polycont >>
rect -20 -145 0 -125
<< locali >>
rect -100 340 -10 350
rect -100 270 -90 340
rect -70 270 -40 340
rect -20 270 -10 340
rect -100 240 -10 270
rect -100 170 -90 240
rect -70 170 -40 240
rect -20 170 -10 240
rect -100 160 -10 170
rect 15 340 55 350
rect 15 270 25 340
rect 45 270 55 340
rect 15 240 55 270
rect 15 170 25 240
rect 45 170 55 240
rect 15 160 55 170
rect 35 95 55 160
rect -100 85 -10 95
rect -100 15 -90 85
rect -70 15 -40 85
rect -20 15 -10 85
rect -100 5 -10 15
rect 15 85 55 95
rect 15 15 25 85
rect 45 15 55 85
rect 15 5 55 15
rect 35 -115 55 5
rect -125 -125 10 -115
rect -125 -135 -20 -125
rect -30 -145 -20 -135
rect 0 -145 10 -125
rect 35 -135 85 -115
rect -30 -155 10 -145
<< viali >>
rect -90 270 -70 340
rect -40 270 -20 340
rect -90 170 -70 240
rect -40 170 -20 240
rect -90 15 -70 85
rect -40 15 -20 85
<< metal1 >>
rect -125 340 85 350
rect -125 270 -90 340
rect -70 270 -40 340
rect -20 270 85 340
rect -125 240 85 270
rect -125 170 -90 240
rect -70 170 -40 240
rect -20 170 85 240
rect -125 160 85 170
rect -125 85 85 95
rect -125 15 -90 85
rect -70 15 -40 85
rect -20 15 85 85
rect -125 -95 85 15
<< labels >>
rlabel metal1 -125 260 -125 260 7 VP
port 3 w
rlabel locali -125 -125 -125 -125 7 A
port 1 w
rlabel locali 85 -125 85 -125 3 Y
port 2 e
rlabel metal1 -125 0 -125 0 7 VN
port 4 w
<< end >>
