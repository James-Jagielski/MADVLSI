magic
tech sky130A
timestamp 1697759168
<< nwell >>
rect -100 360 1835 400
rect -100 -50 1955 360
rect 475 -125 730 -50
rect 1340 -115 1440 -50
rect 640 -130 730 -125
<< nmos >>
rect 85 -560 135 -260
rect 185 -560 235 -260
rect 285 -560 335 -260
rect 385 -560 435 -260
rect 485 -560 535 -260
rect 585 -560 635 -260
rect 685 -560 735 -260
rect 785 -560 835 -260
rect 885 -560 935 -260
rect 985 -560 1035 -260
rect 1085 -560 1135 -260
rect 1185 -560 1235 -260
rect 1285 -560 1335 -260
rect 1385 -560 1435 -260
rect 1485 -560 1535 -260
rect 1585 -560 1635 -260
rect 1685 -560 1735 -260
rect 1785 -560 1835 -260
rect 85 -1085 135 -785
rect 185 -1085 235 -785
rect 285 -1085 335 -785
rect 385 -1085 435 -785
rect 485 -1085 535 -785
rect 585 -1085 635 -785
rect 685 -1085 735 -785
rect 785 -1085 835 -785
rect 885 -1085 935 -785
rect 985 -1085 1035 -785
rect 1085 -1085 1135 -785
rect 1185 -1085 1235 -785
rect 1285 -1085 1335 -785
rect 1385 -1085 1435 -785
rect 1485 -1085 1535 -785
rect 1585 -1085 1635 -785
rect 1685 -1085 1735 -785
rect 1785 -1085 1835 -785
<< pmos >>
rect 85 5 135 305
rect 185 5 235 305
rect 285 5 335 305
rect 385 5 435 305
rect 485 5 535 305
rect 585 5 635 305
rect 685 5 735 305
rect 785 5 835 305
rect 885 5 935 305
rect 985 5 1035 305
rect 1085 5 1135 305
rect 1185 5 1235 305
rect 1285 5 1335 305
rect 1385 5 1435 305
rect 1485 5 1535 305
rect 1585 5 1635 305
rect 1685 5 1735 305
rect 1785 5 1835 305
<< ndiff >>
rect 35 -275 85 -260
rect 35 -545 50 -275
rect 70 -545 85 -275
rect 35 -560 85 -545
rect 135 -275 185 -260
rect 135 -545 150 -275
rect 170 -545 185 -275
rect 135 -560 185 -545
rect 235 -275 285 -260
rect 235 -545 250 -275
rect 270 -545 285 -275
rect 235 -560 285 -545
rect 335 -275 385 -260
rect 335 -545 350 -275
rect 370 -545 385 -275
rect 335 -560 385 -545
rect 435 -275 485 -260
rect 435 -545 450 -275
rect 470 -545 485 -275
rect 435 -560 485 -545
rect 535 -275 585 -260
rect 535 -545 550 -275
rect 570 -545 585 -275
rect 535 -560 585 -545
rect 635 -275 685 -260
rect 635 -545 650 -275
rect 670 -545 685 -275
rect 635 -560 685 -545
rect 735 -275 785 -260
rect 735 -545 750 -275
rect 770 -545 785 -275
rect 735 -560 785 -545
rect 835 -275 885 -260
rect 835 -545 850 -275
rect 870 -545 885 -275
rect 835 -560 885 -545
rect 935 -275 985 -260
rect 935 -545 950 -275
rect 970 -545 985 -275
rect 935 -560 985 -545
rect 1035 -275 1085 -260
rect 1035 -545 1050 -275
rect 1070 -545 1085 -275
rect 1035 -560 1085 -545
rect 1135 -275 1185 -260
rect 1135 -545 1150 -275
rect 1170 -545 1185 -275
rect 1135 -560 1185 -545
rect 1235 -275 1285 -260
rect 1235 -545 1250 -275
rect 1270 -545 1285 -275
rect 1235 -560 1285 -545
rect 1335 -275 1385 -260
rect 1335 -545 1350 -275
rect 1370 -545 1385 -275
rect 1335 -560 1385 -545
rect 1435 -275 1485 -260
rect 1435 -545 1450 -275
rect 1470 -545 1485 -275
rect 1435 -560 1485 -545
rect 1535 -275 1585 -260
rect 1535 -545 1550 -275
rect 1570 -545 1585 -275
rect 1535 -560 1585 -545
rect 1635 -275 1685 -260
rect 1635 -545 1650 -275
rect 1670 -545 1685 -275
rect 1635 -560 1685 -545
rect 1735 -275 1785 -260
rect 1735 -545 1750 -275
rect 1770 -545 1785 -275
rect 1735 -560 1785 -545
rect 1835 -275 1885 -260
rect 1835 -545 1850 -275
rect 1870 -545 1885 -275
rect 1835 -560 1885 -545
rect 35 -800 85 -785
rect 35 -1070 50 -800
rect 70 -1070 85 -800
rect 35 -1085 85 -1070
rect 135 -800 185 -785
rect 135 -1070 150 -800
rect 170 -1070 185 -800
rect 135 -1085 185 -1070
rect 235 -1085 285 -785
rect 335 -800 385 -785
rect 335 -1070 350 -800
rect 370 -1070 385 -800
rect 335 -1085 385 -1070
rect 435 -1085 485 -785
rect 535 -800 585 -785
rect 535 -1070 550 -800
rect 570 -1070 585 -800
rect 535 -1085 585 -1070
rect 635 -1085 685 -785
rect 735 -800 785 -785
rect 735 -1070 750 -800
rect 770 -1070 785 -800
rect 735 -1085 785 -1070
rect 835 -1085 885 -785
rect 935 -800 985 -785
rect 935 -1070 950 -800
rect 970 -1070 985 -800
rect 935 -1085 985 -1070
rect 1035 -1085 1085 -785
rect 1135 -800 1185 -785
rect 1135 -1070 1150 -800
rect 1170 -1070 1185 -800
rect 1135 -1085 1185 -1070
rect 1235 -1085 1285 -785
rect 1335 -800 1385 -785
rect 1335 -1070 1350 -800
rect 1370 -1070 1385 -800
rect 1335 -1085 1385 -1070
rect 1435 -1085 1485 -785
rect 1535 -800 1585 -785
rect 1535 -1070 1550 -800
rect 1570 -1070 1585 -800
rect 1535 -1085 1585 -1070
rect 1635 -1085 1685 -785
rect 1735 -800 1785 -785
rect 1735 -1070 1750 -800
rect 1770 -1070 1785 -800
rect 1735 -1085 1785 -1070
rect 1835 -800 1885 -785
rect 1835 -1070 1850 -800
rect 1870 -1070 1885 -800
rect 1835 -1085 1885 -1070
<< pdiff >>
rect 35 290 85 305
rect 35 20 50 290
rect 70 20 85 290
rect 35 5 85 20
rect 135 290 185 305
rect 135 20 150 290
rect 170 20 185 290
rect 135 5 185 20
rect 235 290 285 305
rect 235 20 250 290
rect 270 20 285 290
rect 235 5 285 20
rect 335 290 385 305
rect 335 20 350 290
rect 370 20 385 290
rect 335 5 385 20
rect 435 290 485 305
rect 435 20 450 290
rect 470 20 485 290
rect 435 5 485 20
rect 535 290 585 305
rect 535 20 550 290
rect 570 20 585 290
rect 535 5 585 20
rect 635 290 685 305
rect 635 20 650 290
rect 670 20 685 290
rect 635 5 685 20
rect 735 290 785 305
rect 735 20 750 290
rect 770 20 785 290
rect 735 5 785 20
rect 835 290 885 305
rect 835 20 850 290
rect 870 20 885 290
rect 835 5 885 20
rect 935 290 985 305
rect 935 20 950 290
rect 970 20 985 290
rect 935 5 985 20
rect 1035 290 1085 305
rect 1035 20 1050 290
rect 1070 20 1085 290
rect 1035 5 1085 20
rect 1135 290 1185 305
rect 1135 20 1150 290
rect 1170 20 1185 290
rect 1135 5 1185 20
rect 1235 290 1285 305
rect 1235 20 1250 290
rect 1270 20 1285 290
rect 1235 5 1285 20
rect 1335 290 1385 305
rect 1335 20 1350 290
rect 1370 20 1385 290
rect 1335 5 1385 20
rect 1435 290 1485 305
rect 1435 20 1450 290
rect 1470 20 1485 290
rect 1435 5 1485 20
rect 1535 290 1585 305
rect 1535 20 1550 290
rect 1570 20 1585 290
rect 1535 5 1585 20
rect 1635 290 1685 305
rect 1635 20 1650 290
rect 1670 20 1685 290
rect 1635 5 1685 20
rect 1735 290 1785 305
rect 1735 20 1750 290
rect 1770 20 1785 290
rect 1735 5 1785 20
rect 1835 295 1885 305
rect 1835 20 1850 295
rect 1870 20 1885 295
rect 1835 5 1885 20
<< ndiffc >>
rect 50 -545 70 -275
rect 150 -545 170 -275
rect 250 -545 270 -275
rect 350 -545 370 -275
rect 450 -545 470 -275
rect 550 -545 570 -275
rect 650 -545 670 -275
rect 750 -545 770 -275
rect 850 -545 870 -275
rect 950 -545 970 -275
rect 1050 -545 1070 -275
rect 1150 -545 1170 -275
rect 1250 -545 1270 -275
rect 1350 -545 1370 -275
rect 1450 -545 1470 -275
rect 1550 -545 1570 -275
rect 1650 -545 1670 -275
rect 1750 -545 1770 -275
rect 1850 -545 1870 -275
rect 50 -1070 70 -800
rect 150 -1070 170 -800
rect 350 -1070 370 -800
rect 550 -1070 570 -800
rect 750 -1070 770 -800
rect 950 -1070 970 -800
rect 1150 -1070 1170 -800
rect 1350 -1070 1370 -800
rect 1550 -1070 1570 -800
rect 1750 -1070 1770 -800
rect 1850 -1070 1870 -800
<< pdiffc >>
rect 50 20 70 290
rect 150 20 170 290
rect 250 20 270 290
rect 350 20 370 290
rect 450 20 470 290
rect 550 20 570 290
rect 650 20 670 290
rect 750 20 770 290
rect 850 20 870 290
rect 950 20 970 290
rect 1050 20 1070 290
rect 1150 20 1170 290
rect 1250 20 1270 290
rect 1350 20 1370 290
rect 1450 20 1470 290
rect 1550 20 1570 290
rect 1650 20 1670 290
rect 1750 20 1770 290
rect 1850 20 1870 295
<< psubdiff >>
rect -15 -275 35 -260
rect -15 -545 0 -275
rect 20 -545 35 -275
rect -15 -560 35 -545
rect 1885 -275 1935 -260
rect 1885 -545 1900 -275
rect 1920 -545 1935 -275
rect 1885 -560 1935 -545
rect -15 -800 35 -785
rect -15 -1070 0 -800
rect 20 -1070 35 -800
rect -15 -1085 35 -1070
rect 1885 -800 1935 -785
rect 1885 -1070 1900 -800
rect 1920 -1070 1935 -800
rect 1885 -1085 1935 -1070
<< nsubdiff >>
rect -15 290 35 305
rect -15 20 0 290
rect 20 20 35 290
rect -15 5 35 20
rect 1885 295 1935 305
rect 1885 20 1900 295
rect 1920 20 1935 295
rect 1885 5 1935 20
<< psubdiffcont >>
rect 0 -545 20 -275
rect 1900 -545 1920 -275
rect 0 -1070 20 -800
rect 1900 -1070 1920 -800
<< nsubdiffcont >>
rect 0 20 20 290
rect 1900 20 1920 295
<< poly >>
rect -20 390 150 400
rect -20 370 -10 390
rect 10 385 150 390
rect 10 370 20 385
rect -20 360 20 370
rect 135 360 150 385
rect 45 350 85 360
rect 45 330 55 350
rect 75 335 85 350
rect 135 345 1635 360
rect 75 330 100 335
rect 45 320 100 330
rect 85 305 135 320
rect 185 305 235 320
rect 285 305 335 345
rect 385 305 435 345
rect 485 305 535 320
rect 585 305 635 320
rect 685 305 735 345
rect 785 305 835 345
rect 885 305 935 320
rect 985 305 1035 320
rect 1085 305 1135 345
rect 1185 305 1235 345
rect 1285 305 1335 320
rect 1385 305 1435 320
rect 1485 305 1535 345
rect 1585 305 1635 345
rect 1840 350 1880 360
rect 1840 335 1850 350
rect 1820 330 1850 335
rect 1870 330 1880 350
rect 1820 320 1880 330
rect 1685 305 1735 320
rect 1785 305 1835 320
rect 85 -10 135 5
rect -10 -20 30 -10
rect -10 -40 0 -20
rect 20 -35 30 -20
rect 185 -35 235 5
rect 285 -10 335 5
rect 385 -10 435 5
rect 485 -35 535 5
rect 585 -35 635 5
rect 685 -10 735 5
rect 785 -10 835 5
rect 885 -35 935 5
rect 985 -35 1035 5
rect 1085 -10 1135 5
rect 1185 -10 1235 5
rect 1285 -35 1335 5
rect 1385 -35 1435 5
rect 1485 -10 1535 5
rect 1585 -10 1635 5
rect 1685 -35 1735 5
rect 1785 -10 1835 5
rect 20 -40 1735 -35
rect -10 -50 1735 -40
rect 2000 -150 2040 -140
rect 2000 -165 2010 -150
rect 105 -170 2010 -165
rect 2030 -170 2040 -150
rect 105 -175 2040 -170
rect 105 -195 115 -175
rect 135 -180 2040 -175
rect 135 -195 145 -180
rect 105 -205 145 -195
rect 40 -215 80 -205
rect 40 -235 50 -215
rect 70 -230 80 -215
rect 70 -235 135 -230
rect 40 -245 135 -235
rect 85 -260 135 -245
rect 185 -260 235 -180
rect 285 -260 335 -245
rect 385 -260 435 -245
rect 485 -260 535 -180
rect 620 -215 660 -205
rect 620 -235 630 -215
rect 650 -235 660 -215
rect 940 -215 980 -205
rect 940 -230 950 -215
rect 620 -245 660 -235
rect 920 -235 950 -230
rect 970 -230 980 -215
rect 1260 -215 1300 -205
rect 970 -235 1000 -230
rect 920 -245 1000 -235
rect 1260 -235 1270 -215
rect 1290 -235 1300 -215
rect 1260 -245 1300 -235
rect 585 -260 635 -245
rect 685 -260 735 -245
rect 785 -260 835 -245
rect 885 -260 935 -245
rect 985 -260 1035 -245
rect 1085 -260 1135 -245
rect 1185 -260 1235 -245
rect 1285 -260 1335 -245
rect 1385 -260 1435 -180
rect 1485 -260 1535 -245
rect 1585 -260 1635 -245
rect 1685 -260 1735 -180
rect 1820 -215 1860 -205
rect 1820 -230 1830 -215
rect 1785 -235 1830 -230
rect 1850 -235 1860 -215
rect 1785 -245 1860 -235
rect 1785 -260 1835 -245
rect 85 -575 135 -560
rect 185 -575 235 -560
rect 25 -675 65 -665
rect 25 -695 35 -675
rect 55 -680 65 -675
rect 285 -680 335 -560
rect 385 -680 435 -560
rect 485 -575 535 -560
rect 585 -575 635 -560
rect 685 -605 735 -560
rect 785 -605 835 -560
rect 885 -575 935 -560
rect 985 -575 1035 -560
rect 1085 -605 1135 -560
rect 1185 -605 1235 -560
rect 1285 -575 1335 -560
rect 1385 -575 1435 -560
rect 485 -615 1235 -605
rect 460 -620 1235 -615
rect 460 -625 500 -620
rect 460 -645 470 -625
rect 490 -645 500 -625
rect 460 -655 500 -645
rect 1485 -680 1535 -560
rect 1585 -680 1635 -560
rect 1685 -575 1735 -560
rect 1785 -575 1835 -560
rect 2000 -665 2040 -655
rect 2000 -680 2010 -665
rect 55 -685 2010 -680
rect 2030 -685 2040 -665
rect 55 -695 2040 -685
rect 25 -705 65 -695
rect 60 -740 100 -730
rect 60 -760 70 -740
rect 90 -760 100 -740
rect 60 -770 100 -760
rect 185 -745 1735 -730
rect 85 -785 135 -770
rect 185 -785 235 -745
rect 285 -785 335 -770
rect 385 -785 435 -770
rect 485 -785 535 -745
rect 585 -785 635 -745
rect 685 -785 735 -770
rect 785 -785 835 -770
rect 885 -785 935 -745
rect 985 -785 1035 -745
rect 1085 -785 1135 -770
rect 1185 -785 1235 -770
rect 1285 -785 1335 -745
rect 1385 -785 1435 -745
rect 1485 -785 1535 -770
rect 1585 -785 1635 -770
rect 1685 -785 1735 -745
rect 1820 -740 1860 -730
rect 1820 -760 1830 -740
rect 1850 -760 1860 -740
rect 1820 -770 1860 -760
rect 1785 -785 1835 -770
rect 85 -1100 135 -1085
rect 185 -1100 235 -1085
rect 15 -1110 55 -1100
rect 15 -1130 25 -1110
rect 45 -1125 55 -1110
rect 205 -1125 220 -1100
rect 285 -1110 335 -1085
rect 385 -1110 435 -1085
rect 485 -1100 535 -1085
rect 585 -1100 635 -1085
rect 285 -1120 435 -1110
rect 285 -1125 350 -1120
rect 45 -1130 220 -1125
rect 15 -1140 220 -1130
rect 340 -1140 350 -1125
rect 370 -1125 435 -1120
rect 685 -1110 735 -1085
rect 785 -1110 835 -1085
rect 885 -1100 935 -1085
rect 985 -1100 1035 -1085
rect 685 -1120 835 -1110
rect 685 -1125 750 -1120
rect 370 -1140 380 -1125
rect 340 -1150 380 -1140
rect 740 -1140 750 -1125
rect 770 -1125 835 -1120
rect 1085 -1110 1135 -1085
rect 1185 -1110 1235 -1085
rect 1285 -1100 1335 -1085
rect 1385 -1100 1435 -1085
rect 1085 -1120 1235 -1110
rect 1085 -1125 1150 -1120
rect 770 -1140 780 -1125
rect 740 -1150 780 -1140
rect 1140 -1140 1150 -1125
rect 1170 -1125 1235 -1120
rect 1485 -1110 1535 -1085
rect 1585 -1110 1635 -1085
rect 1685 -1100 1735 -1085
rect 1785 -1100 1835 -1085
rect 1485 -1120 1635 -1110
rect 1485 -1125 1555 -1120
rect 1170 -1140 1180 -1125
rect 1140 -1150 1180 -1140
rect 1545 -1140 1555 -1125
rect 1575 -1125 1635 -1120
rect 1575 -1140 1585 -1125
rect 1545 -1150 1585 -1140
<< polycont >>
rect -10 370 10 390
rect 55 330 75 350
rect 1850 330 1870 350
rect 0 -40 20 -20
rect 2010 -170 2030 -150
rect 115 -195 135 -175
rect 50 -235 70 -215
rect 630 -235 650 -215
rect 950 -235 970 -215
rect 1270 -235 1290 -215
rect 1830 -235 1850 -215
rect 35 -695 55 -675
rect 470 -645 490 -625
rect 2010 -685 2030 -665
rect 70 -760 90 -740
rect 1830 -760 1850 -740
rect 25 -1130 45 -1110
rect 350 -1140 370 -1120
rect 750 -1140 770 -1120
rect 1150 -1140 1170 -1120
rect 1555 -1140 1575 -1120
<< locali >>
rect -100 390 20 400
rect -100 380 -10 390
rect -20 370 -10 380
rect 10 370 20 390
rect -20 360 20 370
rect 150 380 1770 400
rect 45 350 85 360
rect 45 330 55 350
rect 75 330 85 350
rect 45 320 85 330
rect 50 300 70 320
rect 150 300 170 380
rect 835 350 875 360
rect 835 340 845 350
rect 255 330 845 340
rect 865 330 875 350
rect 255 320 875 330
rect 255 300 275 320
rect 845 300 865 320
rect 950 300 970 380
rect 1045 350 1085 360
rect 1045 330 1055 350
rect 1075 340 1085 350
rect 1075 330 1670 340
rect 1045 320 1670 330
rect 1055 300 1075 320
rect 1650 300 1670 320
rect 1750 300 1770 380
rect 1840 350 1880 360
rect 1840 330 1850 350
rect 1870 330 1880 350
rect 1840 320 1880 330
rect 1860 300 1880 320
rect -10 290 80 300
rect -10 20 0 290
rect 20 20 50 290
rect 70 20 80 290
rect -10 10 80 20
rect 140 290 180 300
rect 140 20 150 290
rect 170 20 180 290
rect 140 10 180 20
rect 240 290 280 300
rect 240 20 250 290
rect 270 20 280 290
rect 240 10 280 20
rect 340 290 380 300
rect 340 20 350 290
rect 370 20 380 290
rect 340 10 380 20
rect 440 290 480 300
rect 440 20 450 290
rect 470 20 480 290
rect 440 10 480 20
rect 540 290 580 300
rect 540 20 550 290
rect 570 20 580 290
rect 540 10 580 20
rect 640 290 680 300
rect 640 20 650 290
rect 670 20 680 290
rect 640 10 680 20
rect 740 290 780 300
rect 740 20 750 290
rect 770 20 780 290
rect 740 10 780 20
rect 840 290 880 300
rect 840 20 850 290
rect 870 20 880 290
rect 840 10 880 20
rect 940 290 980 300
rect 940 20 950 290
rect 970 20 980 290
rect 940 10 980 20
rect 1040 290 1080 300
rect 1040 20 1050 290
rect 1070 20 1080 290
rect 1040 10 1080 20
rect 1140 290 1180 300
rect 1140 20 1150 290
rect 1170 20 1180 290
rect 1140 10 1180 20
rect 1240 290 1280 300
rect 1240 20 1250 290
rect 1270 20 1280 290
rect 1240 10 1280 20
rect 1340 290 1380 300
rect 1340 20 1350 290
rect 1370 20 1380 290
rect 1340 10 1380 20
rect 1440 290 1480 300
rect 1440 20 1450 290
rect 1470 20 1480 290
rect 1440 10 1480 20
rect 1540 290 1580 300
rect 1540 20 1550 290
rect 1570 20 1580 290
rect 1540 10 1580 20
rect 1640 290 1680 300
rect 1640 20 1650 290
rect 1670 20 1680 290
rect 1640 10 1680 20
rect 1740 290 1780 300
rect 1740 20 1750 290
rect 1770 20 1780 290
rect 1740 10 1780 20
rect 1840 295 1930 300
rect 1840 20 1850 295
rect 1870 20 1900 295
rect 1920 20 1930 295
rect 1840 10 1930 20
rect -10 -20 30 -10
rect -10 -30 0 -20
rect -100 -40 0 -30
rect 20 -40 30 -20
rect -100 -50 30 -40
rect 140 -50 160 10
rect 120 -60 160 -50
rect 120 -80 130 -60
rect 150 -80 160 -60
rect 120 -90 160 -80
rect 260 -150 280 10
rect 460 -135 480 10
rect 550 -75 570 10
rect 540 -85 580 -75
rect 540 -105 550 -85
rect 570 -105 580 -85
rect 540 -115 580 -105
rect 640 -135 660 10
rect 840 5 860 10
rect 1260 -135 1280 10
rect 1350 -75 1370 10
rect 1340 -85 1380 -75
rect 1340 -105 1350 -85
rect 1370 -105 1380 -85
rect 1340 -115 1380 -105
rect 1440 -135 1460 10
rect -100 -175 145 -165
rect -100 -185 115 -175
rect 105 -195 115 -185
rect 135 -195 145 -175
rect 105 -205 145 -195
rect 165 -170 280 -150
rect 360 -155 1560 -135
rect 40 -215 80 -205
rect 40 -235 50 -215
rect 70 -235 80 -215
rect 165 -210 185 -170
rect 240 -200 280 -190
rect 240 -210 250 -200
rect 165 -220 250 -210
rect 270 -220 280 -200
rect 165 -225 280 -220
rect 40 -265 80 -235
rect 160 -230 280 -225
rect 160 -245 185 -230
rect 160 -265 180 -245
rect 360 -265 380 -155
rect 540 -200 580 -190
rect 540 -220 550 -200
rect 570 -220 580 -200
rect 540 -230 580 -220
rect 620 -215 660 -205
rect 550 -265 570 -230
rect 620 -235 630 -215
rect 650 -235 660 -215
rect 620 -245 660 -235
rect 940 -215 980 -205
rect 940 -235 950 -215
rect 970 -235 980 -215
rect 940 -245 980 -235
rect 1260 -215 1300 -205
rect 1260 -235 1270 -215
rect 1290 -235 1300 -215
rect 1260 -245 1300 -235
rect 1340 -210 1380 -200
rect 1340 -230 1350 -210
rect 1370 -230 1380 -210
rect 1340 -240 1380 -230
rect 640 -265 660 -245
rect 950 -265 970 -245
rect -10 -275 80 -265
rect -10 -545 0 -275
rect 20 -545 50 -275
rect 70 -545 80 -275
rect -10 -555 80 -545
rect 140 -275 180 -265
rect 140 -545 150 -275
rect 170 -545 180 -275
rect 140 -555 180 -545
rect 240 -275 280 -265
rect 240 -545 250 -275
rect 270 -545 280 -275
rect 240 -555 280 -545
rect 340 -275 380 -265
rect 340 -545 350 -275
rect 370 -545 380 -275
rect 340 -555 380 -545
rect 440 -275 480 -265
rect 440 -545 450 -275
rect 470 -545 480 -275
rect 440 -555 480 -545
rect 540 -275 580 -265
rect 540 -545 550 -275
rect 570 -545 580 -275
rect 540 -555 580 -545
rect 640 -275 680 -265
rect 640 -545 650 -275
rect 670 -545 680 -275
rect 640 -555 680 -545
rect 740 -275 780 -265
rect 740 -545 750 -275
rect 770 -545 780 -275
rect 740 -555 780 -545
rect 840 -275 880 -265
rect 840 -545 850 -275
rect 870 -545 880 -275
rect 840 -555 880 -545
rect 940 -275 980 -265
rect 940 -545 950 -275
rect 970 -545 980 -275
rect 940 -555 980 -545
rect 1040 -275 1080 -260
rect 1260 -265 1280 -245
rect 1350 -265 1370 -240
rect 1540 -265 1560 -155
rect 1650 -150 1670 10
rect 1760 -85 1780 10
rect 1760 -105 1980 -85
rect 1650 -170 1780 -150
rect 1640 -210 1680 -200
rect 1640 -230 1650 -210
rect 1670 -220 1680 -210
rect 1760 -220 1780 -170
rect 1670 -230 1780 -220
rect 1640 -240 1780 -230
rect 1760 -265 1780 -240
rect 1820 -215 1860 -205
rect 1820 -235 1830 -215
rect 1850 -235 1860 -215
rect 1820 -245 1860 -235
rect 1040 -545 1050 -275
rect 1070 -545 1080 -275
rect 1040 -555 1080 -545
rect 1140 -275 1180 -265
rect 1140 -545 1150 -275
rect 1170 -545 1180 -275
rect 1140 -555 1180 -545
rect 1240 -275 1280 -265
rect 1240 -545 1250 -275
rect 1270 -545 1280 -275
rect 1240 -555 1280 -545
rect 1340 -275 1380 -265
rect 1340 -545 1350 -275
rect 1370 -545 1380 -275
rect 1340 -555 1380 -545
rect 1440 -275 1480 -265
rect 1440 -545 1450 -275
rect 1470 -545 1480 -275
rect 1440 -555 1480 -545
rect 1540 -275 1580 -265
rect 1540 -545 1550 -275
rect 1570 -545 1580 -275
rect 1540 -555 1580 -545
rect 1640 -275 1680 -265
rect 1640 -545 1650 -275
rect 1670 -545 1680 -275
rect 1640 -555 1680 -545
rect 1740 -275 1780 -265
rect 1740 -545 1750 -275
rect 1770 -545 1780 -275
rect 1740 -555 1780 -545
rect 1840 -265 1860 -245
rect 1840 -275 1930 -265
rect 1840 -545 1850 -275
rect 1870 -545 1900 -275
rect 1920 -545 1930 -275
rect 1840 -555 1930 -545
rect 260 -575 280 -555
rect 450 -575 470 -555
rect 750 -575 770 -555
rect 1150 -575 1170 -555
rect 1450 -575 1470 -555
rect 1650 -575 1670 -555
rect 260 -595 1670 -575
rect 460 -620 500 -615
rect -100 -625 500 -620
rect -100 -640 470 -625
rect 460 -645 470 -640
rect 490 -645 500 -625
rect 460 -655 500 -645
rect 25 -675 65 -665
rect 1960 -670 1980 -105
rect 2000 -150 2040 -140
rect 2000 -170 2010 -150
rect 2030 -170 2040 -150
rect 2000 -180 2040 -170
rect 25 -685 35 -675
rect -100 -695 35 -685
rect 55 -695 65 -675
rect -100 -705 65 -695
rect 1760 -690 1980 -670
rect 2000 -665 2040 -655
rect 2000 -685 2010 -665
rect 2030 -685 2040 -665
rect 140 -720 180 -710
rect 60 -740 100 -730
rect 60 -760 70 -740
rect 90 -760 100 -740
rect 60 -770 100 -760
rect 140 -740 150 -720
rect 170 -740 180 -720
rect 1320 -715 1360 -705
rect 1320 -725 1330 -715
rect 140 -750 180 -740
rect 560 -735 1330 -725
rect 1350 -735 1360 -715
rect 560 -745 1360 -735
rect 60 -790 80 -770
rect -10 -800 80 -790
rect -10 -1070 0 -800
rect 20 -1070 50 -800
rect 70 -1070 80 -800
rect -10 -1080 80 -1070
rect 140 -790 160 -750
rect 560 -790 580 -745
rect 1340 -790 1360 -745
rect 1760 -790 1780 -690
rect 2000 -695 2040 -685
rect 1820 -740 1860 -730
rect 1820 -760 1830 -740
rect 1850 -760 1860 -740
rect 1820 -770 1860 -760
rect 140 -800 180 -790
rect 140 -1070 150 -800
rect 170 -1070 180 -800
rect 140 -1080 180 -1070
rect 340 -800 380 -790
rect 340 -1070 350 -800
rect 370 -1070 380 -800
rect 340 -1080 380 -1070
rect 540 -800 580 -790
rect 540 -1070 550 -800
rect 570 -1070 580 -800
rect 540 -1080 580 -1070
rect 740 -800 780 -790
rect 740 -1070 750 -800
rect 770 -1070 780 -800
rect 740 -1080 780 -1070
rect 940 -800 980 -790
rect 940 -1070 950 -800
rect 970 -1070 980 -800
rect 940 -1080 980 -1070
rect 1140 -800 1180 -790
rect 1140 -1070 1150 -800
rect 1170 -1070 1180 -800
rect 1140 -1080 1180 -1070
rect 1340 -800 1380 -790
rect 1340 -1070 1350 -800
rect 1370 -1070 1380 -800
rect 1340 -1080 1380 -1070
rect 1540 -800 1580 -790
rect 1540 -1070 1550 -800
rect 1570 -1070 1580 -800
rect 1540 -1080 1580 -1070
rect 1740 -800 1780 -790
rect 1740 -1070 1750 -800
rect 1770 -1070 1780 -800
rect 1740 -1080 1780 -1070
rect 1840 -790 1860 -770
rect 1840 -800 1930 -790
rect 1840 -1070 1850 -800
rect 1870 -1070 1900 -800
rect 1920 -1070 1930 -800
rect 1840 -1080 1930 -1070
rect 15 -1110 55 -1100
rect -100 -1140 -15 -1120
rect 15 -1130 25 -1110
rect 45 -1130 55 -1110
rect 15 -1140 55 -1130
rect 160 -1120 180 -1080
rect 340 -1120 380 -1110
rect 740 -1120 780 -1110
rect 945 -1120 975 -1080
rect 1140 -1120 1180 -1110
rect 1545 -1120 1585 -1110
rect 1745 -1120 1765 -1080
rect 160 -1140 350 -1120
rect 370 -1140 750 -1120
rect 770 -1140 1150 -1120
rect 1170 -1140 1555 -1120
rect 1575 -1140 1765 -1120
rect 340 -1150 380 -1140
rect 740 -1150 780 -1140
rect 1140 -1150 1180 -1140
rect 1545 -1150 1585 -1140
<< viali >>
rect 845 330 865 350
rect 1055 330 1075 350
rect 0 20 20 290
rect 50 20 70 290
rect 350 20 370 290
rect 750 20 770 290
rect 1150 20 1170 290
rect 1550 20 1570 290
rect 1850 20 1870 295
rect 1900 20 1920 295
rect 130 -80 150 -60
rect 550 -105 570 -85
rect 1350 -105 1370 -85
rect 250 -220 270 -200
rect 550 -220 570 -200
rect 1350 -230 1370 -210
rect 0 -545 20 -275
rect 50 -545 70 -275
rect 650 -545 670 -275
rect 850 -545 870 -275
rect 950 -545 970 -275
rect 1650 -230 1670 -210
rect 1050 -545 1070 -275
rect 1250 -545 1270 -275
rect 1850 -545 1870 -275
rect 1900 -545 1920 -275
rect 150 -740 170 -720
rect 1330 -735 1350 -715
rect 0 -1070 20 -800
rect 50 -1070 70 -800
rect 350 -1070 370 -800
rect 750 -1070 770 -800
rect 1150 -1070 1170 -800
rect 1550 -1070 1570 -800
rect 1850 -1070 1870 -800
rect 1900 -1070 1920 -800
<< metal1 >>
rect 835 350 1085 360
rect 835 330 845 350
rect 865 340 1055 350
rect 865 330 875 340
rect 835 320 875 330
rect 1045 330 1055 340
rect 1075 330 1085 350
rect 1045 320 1085 330
rect -100 295 1935 305
rect -100 290 1850 295
rect -100 20 0 290
rect 20 20 50 290
rect 70 20 350 290
rect 370 20 750 290
rect 770 20 1150 290
rect 1170 20 1550 290
rect 1570 20 1850 290
rect 1870 20 1900 295
rect 1920 20 1935 295
rect -100 5 1935 20
rect 120 -60 160 -50
rect 120 -70 130 -60
rect -65 -80 130 -70
rect 150 -80 160 -60
rect -65 -90 160 -80
rect 540 -85 1995 -75
rect -65 -640 -45 -90
rect 540 -105 550 -85
rect 570 -105 1350 -85
rect 1370 -105 1995 -85
rect 540 -115 1995 -105
rect 240 -200 280 -190
rect 240 -220 250 -200
rect 270 -210 280 -200
rect 540 -200 580 -190
rect 540 -210 550 -200
rect 270 -220 550 -210
rect 570 -220 580 -200
rect 240 -230 580 -220
rect 1340 -210 1680 -200
rect 1340 -230 1350 -210
rect 1370 -230 1650 -210
rect 1670 -230 1680 -210
rect 1340 -240 1680 -230
rect 1895 -260 1945 -255
rect -30 -275 1945 -260
rect -30 -545 0 -275
rect 20 -545 50 -275
rect 70 -545 650 -275
rect 670 -545 850 -275
rect 870 -545 950 -275
rect 970 -545 1050 -275
rect 1070 -545 1250 -275
rect 1270 -545 1850 -275
rect 1870 -545 1900 -275
rect 1920 -545 1945 -275
rect -30 -560 1945 -545
rect -30 -565 20 -560
rect -65 -665 165 -640
rect 140 -710 165 -665
rect 140 -720 180 -710
rect 140 -740 150 -720
rect 170 -740 180 -720
rect 140 -750 180 -740
rect 235 -785 1285 -560
rect 1960 -660 1995 -115
rect 1320 -690 1995 -660
rect 1320 -715 1360 -690
rect 1320 -735 1330 -715
rect 1350 -735 1360 -715
rect 1320 -745 1360 -735
rect -100 -800 1935 -785
rect -100 -1070 0 -800
rect 20 -1070 50 -800
rect 70 -1070 350 -800
rect 370 -1070 750 -800
rect 770 -1070 1150 -800
rect 1170 -1070 1550 -800
rect 1570 -1070 1850 -800
rect 1870 -1070 1900 -800
rect 1920 -1070 1935 -800
rect -100 -1085 1935 -1070
<< labels >>
rlabel locali -100 390 -100 390 7 Vbp
port 1 w
rlabel locali -100 -40 -100 -40 7 Vcp
port 3 w
rlabel locali -100 -175 -100 -175 7 V1
port 4 w
rlabel locali -100 -630 -100 -630 7 Vbn
port 5 w
rlabel locali -100 -695 -100 -695 7 V2
port 6 w
rlabel metal1 -100 -935 -100 -935 7 GND
port 7 w
rlabel locali -100 -1130 -100 -1130 7 Vcn
port 8 w
rlabel metal1 -100 160 -100 160 7 VDD
port 2 w
rlabel metal1 1995 -410 1995 -410 3 Vout
port 9 e
<< end >>
