* NGSPICE file created from Cascode_voltage_bias.ext - technology: sky130A


X0 a_2640_2790# a_2640_2790# Vcp VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X1 Vcp a_2140_2820# a_2140_2820# VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X2 Vcp a_2640_2790# VDD VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X3 a_2690_4480# Vbp a_2540_4480# VDD sky130_fd_pr__pfet_01v8 ad=0.75 pd=6.25 as=0.75 ps=6.25 w=6 l=0.5
X4 a_2840_4480# Vbp a_2690_4480# VDD sky130_fd_pr__pfet_01v8 ad=0.75 pd=6.25 as=0.75 ps=6.25 w=6 l=0.5
X5 a_3240_1290# Vbn a_3090_1290# GND sky130_fd_pr__nfet_01v8 ad=0.75 pd=6.25 as=0.75 ps=6.25 w=6 l=0.5
X6 VDD Vbp Vcn VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X7 a_3890_1290# Vbn a_3740_1290# GND sky130_fd_pr__nfet_01v8 ad=0.75 pd=6.25 as=0.75 ps=6.25 w=6 l=0.5
X8 a_4040_1290# Vbn a_3890_1290# GND sky130_fd_pr__nfet_01v8 ad=0.75 pd=6.25 as=0.75 ps=6.25 w=6 l=0.5
X9 GND GND Vbn GND sky130_fd_pr__nfet_01v8 ad=3 pd=13 as=1.5 ps=6.5 w=6 l=0.5
X10 Vbp VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=3 ps=13 w=6 l=0.5
X11 Vbn Vbp VDD VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X12 VDD Vbp Vbn VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X13 a_2140_2820# Vbn GND GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X14 a_2340_n260# a_2640_n290# a_2640_n290# GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X15 Vcn Vbp VDD VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X16 a_2640_1290# Vbn GND GND sky130_fd_pr__nfet_01v8 ad=0.75 pd=6.25 as=1.5 ps=6.5 w=6 l=0.5
X17 a_2340_n260# GND GND GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X18 a_3190_4480# Vbp a_2640_n290# VDD sky130_fd_pr__pfet_01v8 ad=0.75 pd=6.25 as=1.5 ps=6.5 w=6 l=0.5
X19 a_3340_4480# Vbp a_3190_4480# VDD sky130_fd_pr__pfet_01v8 ad=0.75 pd=6.25 as=0.75 ps=6.25 w=6 l=0.5
X20 VDD VDD a_2140_2820# VDD sky130_fd_pr__pfet_01v8 ad=3 pd=13 as=1.5 ps=6.5 w=6 l=0.5
X21 a_2140_2820# GND GND GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X22 a_2640_n290# a_2640_n290# a_2340_n260# GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X23 Vbn Vbn GND GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X24 a_2640_n290# a_2640_n290# a_2340_n260# GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X25 a_2640_2790# a_2640_2790# Vcp VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X26 VDD a_2640_2790# Vcp VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X27 GND Vbn Vbn GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X28 a_2140_2820# a_2140_2820# Vcp VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X29 a_2640_2790# Vbn a_3240_1290# GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=0.75 ps=6.25 w=6 l=0.5
X30 a_2340_n260# Vcn Vcn GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X31 a_2640_n290# Vbp a_2840_4480# VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=0.75 ps=6.25 w=6 l=0.5
X32 Vcp a_2640_2790# a_2640_2790# VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X33 a_2340_n260# a_2640_n290# GND GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X34 Vcp a_2640_2790# a_2640_2790# VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X35 Vcp a_2640_2790# a_2640_2790# VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X36 a_2140_2820# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=3 ps=13 w=6 l=0.5
X37 a_2790_1290# Vbn a_2640_1290# GND sky130_fd_pr__nfet_01v8 ad=0.75 pd=6.25 as=0.75 ps=6.25 w=6 l=0.5
X38 a_2940_1290# Vbn a_2790_1290# GND sky130_fd_pr__nfet_01v8 ad=0.75 pd=6.25 as=0.75 ps=6.25 w=6 l=0.5
X39 a_3490_4480# Vbp a_3340_4480# VDD sky130_fd_pr__pfet_01v8 ad=0.75 pd=6.25 as=0.75 ps=6.25 w=6 l=0.5
X40 a_3640_4480# Vbp a_3490_4480# VDD sky130_fd_pr__pfet_01v8 ad=0.75 pd=6.25 as=0.75 ps=6.25 w=6 l=0.5
X41 VDD VDD Vcp VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X42 VDD VDD Vbp VDD sky130_fd_pr__pfet_01v8 ad=3 pd=13 as=1.5 ps=6.5 w=6 l=0.5
X43 a_2640_2790# a_2640_2790# Vcp VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X44 a_2240_4480# Vbp VDD VDD sky130_fd_pr__pfet_01v8 ad=0.75 pd=6.25 as=1.5 ps=6.5 w=6 l=0.5
X45 GND GND Vcn GND sky130_fd_pr__nfet_01v8 ad=3 pd=13 as=1.5 ps=6.5 w=6 l=0.5
X46 Vcn VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X47 VDD Vbp Vbp VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X48 Vbn VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X49 a_2640_n290# a_2640_n290# a_2340_n260# GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X50 VDD VDD Vbn VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X51 Vbp Vbp VDD VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X52 GND GND a_2140_2820# GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X53 GND a_2640_n290# a_2340_n260# GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X54 VDD VDD Vcn VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X55 a_3090_1290# Vbn a_2940_1290# GND sky130_fd_pr__nfet_01v8 ad=0.75 pd=6.25 as=0.75 ps=6.25 w=6 l=0.5
X56 Vcn Vcn a_2340_n260# GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X57 a_3790_4480# Vbp a_3640_4480# VDD sky130_fd_pr__pfet_01v8 ad=0.75 pd=6.25 as=0.75 ps=6.25 w=6 l=0.5
X58 a_4190_1290# Vbn a_4040_1290# GND sky130_fd_pr__nfet_01v8 ad=0.75 pd=6.25 as=0.75 ps=6.25 w=6 l=0.5
X59 GND Vbn a_4190_1290# GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=0.75 ps=6.25 w=6 l=0.5
X60 a_2340_n260# a_2640_n290# a_2640_n290# GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X61 VDD Vbp a_3790_4480# VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=0.75 ps=6.25 w=6 l=0.5
X62 GND Vbn a_2140_2820# GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X63 a_2340_n260# a_2640_n290# a_2640_n290# GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X64 a_2390_4480# Vbp a_2240_4480# VDD sky130_fd_pr__pfet_01v8 ad=0.75 pd=6.25 as=0.75 ps=6.25 w=6 l=0.5
X65 Vcp a_2640_2790# a_2640_2790# VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X66 Vbn GND GND GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=3 ps=13 w=6 l=0.5
X67 a_2340_n260# a_2640_n290# a_2640_n290# GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X68 a_2540_4480# Vbp a_2390_4480# VDD sky130_fd_pr__pfet_01v8 ad=0.75 pd=6.25 as=0.75 ps=6.25 w=6 l=0.5
X69 Vcp VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X70 a_3590_1290# Vbn a_2640_2790# GND sky130_fd_pr__nfet_01v8 ad=0.75 pd=6.25 as=1.5 ps=6.5 w=6 l=0.5
X71 Vcn GND GND GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=3 ps=13 w=6 l=0.5
X72 a_3740_1290# Vbn a_3590_1290# GND sky130_fd_pr__nfet_01v8 ad=0.75 pd=6.25 as=0.75 ps=6.25 w=6 l=0.5
X73 GND GND a_2340_n260# GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X74 a_2640_2790# a_2640_2790# Vcp VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X75 a_2640_n290# a_2640_n290# a_2340_n260# GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
.ends

