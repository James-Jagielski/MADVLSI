* NGSPICE file created from AND2.ext - technology: sky130A

.subckt inverter A Y VP VN
X0 Y A VP VP sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X1 Y A VN VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
.ends

.subckt NAND A B Y VP VN
X0 Y A VP VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=1 ps=5 w=2 l=0.15
X1 VP B Y VP sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=0.5 ps=2.5 w=2 l=0.15
X2 Y B a_80_n200# VN sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0.25 ps=2.25 w=2 l=0.15
X3 a_80_n200# A VN VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=2.25 as=1 ps=5 w=2 l=0.15
.ends


* Top level circuit AND2

Xinverter_0 NAND_0/Y inverter_0/Y NAND_0/VP VSUBS inverter
XNAND_0 NAND_0/A NAND_0/B NAND_0/Y NAND_0/VP VSUBS NAND
.end

