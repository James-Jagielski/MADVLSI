magic
tech sky130A
timestamp 1694482200
<< nwell >>
rect -125 135 150 375
<< nmos >>
rect 25 -100 40 100
rect 65 -100 80 100
<< pmos >>
rect 0 155 15 355
rect 65 155 80 355
<< ndiff >>
rect -25 85 25 100
rect -25 15 -10 85
rect 10 15 25 85
rect -25 -15 25 15
rect -25 -85 -10 -15
rect 10 -85 25 -15
rect -25 -100 25 -85
rect 40 -100 65 100
rect 80 85 130 100
rect 80 15 95 85
rect 115 15 130 85
rect 80 -15 130 15
rect 80 -85 95 -15
rect 115 -85 130 -15
rect 80 -100 130 -85
<< pdiff >>
rect -50 340 0 355
rect -50 270 -35 340
rect -15 270 0 340
rect -50 240 0 270
rect -50 170 -35 240
rect -15 170 0 240
rect -50 155 0 170
rect 15 340 65 355
rect 15 270 30 340
rect 50 270 65 340
rect 15 240 65 270
rect 15 170 30 240
rect 50 170 65 240
rect 15 155 65 170
rect 80 340 130 355
rect 80 270 95 340
rect 115 270 130 340
rect 80 240 130 270
rect 80 170 95 240
rect 115 170 130 240
rect 80 155 130 170
<< ndiffc >>
rect -10 15 10 85
rect -10 -85 10 -15
rect 95 15 115 85
rect 95 -85 115 -15
<< pdiffc >>
rect -35 270 -15 340
rect -35 170 -15 240
rect 30 270 50 340
rect 30 170 50 240
rect 95 270 115 340
rect 95 170 115 240
<< psubdiff >>
rect -75 85 -25 100
rect -75 15 -60 85
rect -40 15 -25 85
rect -75 -15 -25 15
rect -75 -85 -60 -15
rect -40 -85 -25 -15
rect -75 -100 -25 -85
<< nsubdiff >>
rect -100 340 -50 355
rect -100 270 -85 340
rect -65 270 -50 340
rect -100 240 -50 270
rect -100 170 -85 240
rect -65 170 -50 240
rect -100 155 -50 170
<< psubdiffcont >>
rect -60 15 -40 85
rect -60 -85 -40 -15
<< nsubdiffcont >>
rect -85 270 -65 340
rect -85 170 -65 240
<< poly >>
rect 0 355 15 370
rect 65 355 80 370
rect 0 125 15 155
rect 0 110 40 125
rect 25 100 40 110
rect 65 100 80 155
rect 25 -115 40 -100
rect 0 -125 40 -115
rect 0 -145 10 -125
rect 30 -145 40 -125
rect 0 -155 40 -145
rect 65 -180 80 -100
rect 40 -190 80 -180
rect 40 -210 50 -190
rect 70 -210 80 -190
rect 40 -220 80 -210
<< polycont >>
rect 10 -145 30 -125
rect 50 -210 70 -190
<< locali >>
rect -95 340 -5 350
rect -95 270 -85 340
rect -65 270 -35 340
rect -15 270 -5 340
rect -95 240 -5 270
rect -95 170 -85 240
rect -65 170 -35 240
rect -15 170 -5 240
rect -95 160 -5 170
rect 20 340 60 350
rect 20 270 30 340
rect 50 270 60 340
rect 20 240 60 270
rect 20 170 30 240
rect 50 170 60 240
rect 20 160 60 170
rect 85 340 125 350
rect 85 270 95 340
rect 115 270 125 340
rect 85 240 125 270
rect 85 170 95 240
rect 115 170 125 240
rect 85 160 125 170
rect 40 95 60 160
rect -70 85 20 95
rect -70 15 -60 85
rect -40 15 -10 85
rect 10 15 20 85
rect 40 85 125 95
rect 40 75 95 85
rect -70 -15 20 15
rect -70 -85 -60 -15
rect -40 -85 -10 -15
rect 10 -85 20 -15
rect -70 -95 20 -85
rect 85 15 95 75
rect 115 15 125 85
rect 85 -15 125 15
rect 85 -85 95 -15
rect 115 -85 125 -15
rect 85 -95 125 -85
rect 105 -115 125 -95
rect -125 -125 40 -115
rect -125 -135 10 -125
rect 0 -145 10 -135
rect 30 -145 40 -125
rect 105 -135 150 -115
rect 0 -155 40 -145
rect -125 -190 80 -180
rect -125 -200 50 -190
rect 40 -210 50 -200
rect 70 -210 80 -190
rect 40 -220 80 -210
<< viali >>
rect -85 270 -65 340
rect -35 270 -15 340
rect -85 170 -65 240
rect -35 170 -15 240
rect 95 270 115 340
rect 95 170 115 240
rect -60 15 -40 85
rect -10 15 10 85
rect -60 -85 -40 -15
rect -10 -85 10 -15
<< metal1 >>
rect -125 340 150 350
rect -125 270 -85 340
rect -65 270 -35 340
rect -15 270 95 340
rect 115 270 150 340
rect -125 240 150 270
rect -125 170 -85 240
rect -65 170 -35 240
rect -15 170 95 240
rect 115 170 150 240
rect -125 160 150 170
rect -125 85 150 95
rect -125 15 -60 85
rect -40 15 -10 85
rect 10 15 150 85
rect -125 -15 150 15
rect -125 -85 -60 -15
rect -40 -85 -10 -15
rect 10 -85 150 -15
rect -125 -95 150 -85
<< labels >>
rlabel locali -125 -125 -125 -125 7 A
port 1 w
rlabel locali -125 -190 -125 -190 7 B
port 2 w
rlabel locali 150 -125 150 -125 3 Y
port 3 e
rlabel metal1 -125 255 -125 255 7 VP
port 4 w
rlabel metal1 -125 0 -125 0 7 VN
port 5 w
<< end >>
